netcdf NCEI_TimeSeries_Orthogonal {
dimensions:
       time = 1;
variables:
        double time(time) ;
                time:long_name = "Time" ; 
                time:standard_name = "time" ; 
                time:units = "seconds since 1970-01-01 00:00:00 0:00" ; 
                time:calendar = "gregorian" ; 
                time:axis = "T" ; 
                time:ancillary_variables = "" ; 
                time:comment = "Time" ; 
        float lat ;
                lat:long_name = "Latitude" ; 
                lat:standard_name = "latitude" ; 
                lat:units = "degrees_north" ; 
                lat:axis = "Y" ; 
                lat:valid_min = -90.0f ; 
                lat:valid_max = 90.0f ; 
                lat:_FillValue = -9999.0f;
                lat:ancillary_variables = "" ; 
                lat:comment = "" ; 
       float lon ; 
                lon:long_name = "Longitude" ; 
                lon:standard_name = "longitude" ; 
                lon:units = "degrees_east" ; 
                lon:axis = "X" ; 
                lon:valid_min = -180.0f ; 
                lon:valid_max = 180.0f ; 
                lon:_FillValue = -9999.0f;
                lon:ancillary_variables = "" ; 
                lon:comment = "" ; 
        float z ;
                z:long_name = "Depth Below Sea Surface" ; 
                z:standard_name = "depth" ; 
                z:units = "m" ; 
                z:axis = "Z" ; 
                z:positive = "down" ; 
                z:valid_min = 0.0f ; 
                z:valid_max = 1000.0f ; 
                z:_FillValue = -9999.0f;
                z:ancillary_variables = "" ; 
                z:comment = "" ; 

        float temperature(time) ;
                temperature:long_name = "Sea Water Temperature" ; 
                temperature:standard_name = "sea_water_temperature" ; 
                temperature:ncei_name = "" ; 
                temperature:units = "" ; 
                temperature:scale_factor = 0.0f ; 
                temperature:add_offset = 0.0f ; 
                temperature:_FillValue = 0.0f ; 
                temperature:missing_value = 0.0f ; 
                temperature:valid_min = 0.0f ; 
                temperature:valid_max = 0.0f ; 
                temperature:coordinates = "time lat lon z" ; 
                temperature:coverage_content_type = "" ; 
                temperature:grid_mapping = "crs" ; 
                temperature:source = "" ; 
                temperature:references = "" ; 
                temperature: cell_methods = "" ; 
                temperature:ancillary_variables = "temperature_qc" ; 
                temperature:platform = "platform_id" ; 
                temperature:instrument = "instrument_id";
                temperature:comment = "" ; 

        int temperature_qc(time);  
                temperature_qc:standard_name= "" ; 
                temperature_qc:long_name = "" ; 
                temperature_qc:flag_values = ""; 
                temperature_qc:flag_meanings = "" ; 
                temperature_qc:references = "" ; 
                temperature_qc:comment = "" ; 

        int platform_id; 
                platform_id:long_name = "" ; 
                platform_id:comment = "" ; 
                platform_id:call_sign = "" ; 
                platform_id:ncei_code = ""; 
                platform_id:wmo_code = "";
                platform_id:imo_code  = "";

        int instrument_id; 
                instrument_id:long_name = "" ; 
                instrument_id:comment = "" ; 
        double crs; 
                crs:grid_mapping_name = "latitude_longitude"; 
                crs:epsg_code = "EPSG:4326" ; 
                crs:semi_major_axis = 6378137.0d ; 
                crs:inverse_flattening = 298.257223563d ; 



        :ncei_template_version = "NCEI_NetCDF_TimeSeries_Orthogonal_Template_v2.0" ; 
        :featureType = "timeSeries" ; 
        :title = "" ; 
        :summary = "" ; 
        :keywords = "" ; 
        :Conventions = "CF-1.6, ACDD-1.3" ; 
        :id = "" ; 
       :naming_authority = "" ; 
       :history = "" ; 
       :source = "" ; 
       :processing_level = "" ; 
       :comment = "" ; 
       :acknowledgment = "" ; 
       :license = "" ; 
       :standard_name_vocabulary = "CF Standard Name Table vNN" ; 
       :date_created = "" ; 
       :creator_name = "" ; 
       :creator_email = "" ; 
       :creator_url = "" ; 
       :institution = "" ; 
       :project = "" ; 
       :publisher_name = "" ; 
       :publisher_email = "" ; 
       :publisher_url = "" ; 
       :geospatial_bounds = "" ; 
       :geospatial_bounds_crs = "" ; 
       :geospatial_bounds_vertical_crs = "" ; 
       :geospatial_lat_min = 0.0d ; 
       :geospatial_lat_max = 0.0d ; 
       :geospatial_lon_min = 0.0d ; 
       :geospatial_lon_max = 0.0d ; 
       :geospatial_vertical_min = 0.0d ; 
       :geospatial_vertical_max = 0.0d ; 
       :geospatial_vertical_positive = "" ; 
       :time_coverage_start = "" ; 
       :time_coverage_end = "" ; 
       :time_coverage_duration = "" ; 
       :time_coverage_resolution = "" ; 
       :uuid = "" ; 
       :sea_name = "" ; 
       :creator_type = "" ; 
       :creator_institution = "" ; 
       :publisher_type = "" ; 
       :publisher_institution = "" ; 
       :program = "" ; 
       :contributor_name = "" ; 
       :contributor_role = "" ; 
       :geospatial_lat_units = "degrees_north" ; 
       :geospatial_lon_units = "degrees_east"; 
       :geospatial_vertical_units = "" ; 
       :date_modified = "" ; 
       :date_issued = "" ; 
       :date_metadata_modified = "" ; 
       :product_version = "" ; 
       :keywords_vocabulary = "" ; 
       :platform = "" ; 
       :platform_vocabulary = "" ; 
       :instrument = "" ; 
       :instrument_vocabulary = "" ; 
       :cdm_data_type = "Station" ; 
       :metadata_link = "" ; 
       :references = "" ; 
       
      
}

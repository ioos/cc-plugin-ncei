netcdf usgs_internal_wave_timeSeries {
dimensions:
	time = 38990 ;
	nzMax = 5 ;
	station = 1 ;
variables:
	int station(station) ;
		station:long_name = "" ;
		station:cf_role = "timeseries_id" ;
	double time(time) ;
		time:long_name = "time [seconds since 1970 00:00:00 00:00]" ;
		time:standard_name = "time" ;
		time:units = "seconds since 1970-01-01 00:00:00 00:00" ;
		time:calendar = "gregorian" ;
		time:axis = "T" ;
		time:type = "EVEN" ;
		time:epic_code = 624. ;
		time:comment = " " ;
		time:ancillary_variables = " " ;
	double z(station, time, nzMax) ;
		z:long_name = "Depth [m]" ;
		z:standard_name = "depth" ;
		z:units = "m" ;
		z:axis = "Z" ;
		z:positive = "down" ;
		z:valid_min = 0.f ;
		z:valid_max = 15000.f ;
		z:ancillary_variables = "instrument_1" ;
		z:type = "EVEN" ;
		z:epic_code = 3. ;
		z:comment = "" ;
	double lon(station) ;
		lon:long_name = "longitude [degrees east]" ;
		lon:standard_name = "longitude" ;
		lon:units = "degrees_east" ;
		lon:axis = "X" ;
		lon:valid_min = -180.f ;
		lon:valid_max = 180.f ;
		lon:ancillary_variables = "instrument_2" ;
		lon:type = "EVEN" ;
		lon:epic_code = 502. ;
		lon:comment = "" ;
	double lat(station) ;
		lat:long_name = "latitude [degrees north]" ;
		lat:standard_name = "latitude" ;
		lat:units = "degrees_north" ;
		lat:axis = "Y" ;
		lat:valid_min = -90.f ;
		lat:valid_max = 90.f ;
		lat:ancillary_variables = "instrument_2" ;
		lat:type = "EVEN" ;
		lat:epic_code = 500. ;
		lat:comment = "" ;
	double T_20(station, time, nzMax) ;
		T_20:long_name = "TEMPERATURE (C)" ;
		T_20:standard_name = "sea_water_temperature" ;
		T_20:nodc_name = "TEMPERATURE" ;
		T_20:units = "Celsius" ;
		T_20:scale_factor = 1.f ;
		T_20:add_offset = 0.f ;
		T_20:_FillValue = NaN ;
		T_20:valid_min = 0. ;
		T_20:valid_max = 100. ;
		T_20:data_min = 6.98519992828369 ;
		T_20:data_max = 18.1453990936279 ;
		T_20:coordinates = "time lon lat z" ;
		T_20:grid_mapping = "crs" ;
		T_20:source = "" ;
		T_20:references = "http://www.nodc.noaa.gov/archive/arc0033/0061443/1.1/" ;
		T_20:cell_methods = "time: point longitude: point latitude: point z: point" ;
		T_20:ancillary_variables = "instrument_1" ;
		T_20:type = "" ;
		T_20:epic_code = 20. ;
		T_20:comment = "Data were reformatted from original EPIC conventions NetCDF data" ;
	double C_51(station, time, nzMax) ;
		C_51:long_name = "CONDUCTIVITY             " ;
		C_51:standard_name = "sea_water_electrical_conductivity" ;
		C_51:nodc_name = "CONDUCTIVITY" ;
		C_51:units = "S/m" ;
		C_51:scale_factor = 1.f ;
		C_51:add_offset = 0.f ;
		C_51:_FillValue = NaN ;
		C_51:valid_min = 0. ;
		C_51:valid_max = 10. ;
		C_51:data_min = 3.20242595672607 ;
		C_51:data_max = 4.08073616027832 ;
		C_51:coordinates = "time lat lon z" ;
		C_51:grid_mapping = "crs" ;
		C_51:source = "" ;
		C_51:references = "http://www.nodc.noaa.gov/archive/arc0033/0061443/1.1/" ;
		C_51:cell_methods = "time: point longitude: point latitude: point z: point" ;
		C_51:ancillary_variables = "instrument_1" ;
		C_51:type = "" ;
		C_51:epic_code = 51. ;
		C_51:comment = "Data were reformatted from original EPIC conventions NetCDF data" ;
	double S_40(station, time, nzMax) ;
		S_40:long_name = "SALINITY (PPT)           " ;
		S_40:standard_name = "sea_water_salinity" ;
		S_40:nodc_name = "SALINITY" ;
		S_40:units = "0.001" ;
		S_40:scale_factor = 1.f ;
		S_40:add_offset = 0.f ;
		S_40:_FillValue = NaN ;
		S_40:valid_min = 0. ;
		S_40:valid_max = 40. ;
		S_40:data_min = 28.3021602630615 ;
		S_40:data_max = 33.0736122131348 ;
		S_40:coordinates = "time lat lon z" ;
		S_40:grid_mapping = "crs" ;
		S_40:source = "" ;
		S_40:references = "http://www.nodc.noaa.gov/archive/arc0033/0061443/1.1/" ;
		S_40:cell_methods = "time: point longitude: point latitude: point z: point" ;
		S_40:ancillary_variables = "instrument_1" ;
		S_40:type = "" ;
		S_40:epic_code = 40. ;
		S_40:comment = "Data were reformatted from original EPIC conventions NetCDF data" ;
	double STH_71(station, time, nzMax) ;
		STH_71:long_name = "SIGMA-THETA (KG/M**3)    " ;
		STH_71:standard_name = "sea_water_sigma_theta" ;
		STH_71:nodc_name = "SIGMA-THETA" ;
		STH_71:units = "kg m-3" ;
		STH_71:scale_factor = 1.f ;
		STH_71:add_offset = 0.f ;
		STH_71:_FillValue = NaN ;
		STH_71:valid_min = 0. ;
		STH_71:valid_max = 40. ;
		STH_71:data_min = 20.5344085693359 ;
		STH_71:data_max = 25.1763973236084 ;
		STH_71:coordinates = "time lat lon z" ;
		STH_71:grid_mapping = "crs" ;
		STH_71:source = "" ;
		STH_71:references = "http://www.nodc.noaa.gov/archive/arc0033/0061443/1.1/" ;
		STH_71:cell_methods = "time: point longitude: point latitude: point z: point" ;
		STH_71:ancillary_variables = "instrument_1" ;
		STH_71:type = "" ;
		STH_71:epic_code = 71. ;
		STH_71:comment = "Data were reformatted from original EPIC conventions NetCDF data" ;
	int instrument_1(station) ;
		instrument_1:long_name = "Seabird SBE16 Seacat serial number" ;
		instrument_1:nodc_name = "CTD - specific model" ;
		instrument_1:make_model = "Seabird SBE16 Seacat" ;
		instrument_1:calibration_date = "" ;
		instrument_1:comment = "" ;
	int instrument_2(station) ;
		instrument_2:long_name = "Global Positioning System" ;
		instrument_2:nodc_name = "GPS" ;
		instrument_2:make_model = "" ;
		instrument_2:serial_number = "" ;
		instrument_2:calibration_date = "" ;
		instrument_2:comment = "" ;
	int platform ;
		platform:long_name = "usgs mooring 5391" ;
		platform:comment = "usgs mooring" ;
		platform:call_sign = "" ;
		platform:nodc_code = "" ;
		platform:wmo_code = "" ;
		platform:imo_code = "" ;
	int crs ;
		crs:grid_mapping_name = "latitude_longitude" ;
		crs:longitude_of_prime_meridian = 0. ;
		crs:epsg_code = "EPSG:4326" ;
		crs:semi_major_axis = 6378137. ;
		crs:inverse_flattening = 298.257223563 ;

// global attributes:
		:Conventions = "CF-1.6" ;
		:Metadata_Conventions = "Unidata Dataset Discovery v1.0" ;
		:featureType = "timeSeriesProfile" ;
		:cdm_data_type = "Station" ;
		:nodc_template_version = "NODC_NetCDF_TimeSeriesProfile_IncompleteVertical_OrthogonalTemporal_Template_v1.1" ;
		:standard_name_vocabulary = "NetCDF Climate and Forecast (CF) Metadata Convention Standard Name Table v23" ;
		:title = "Temperature and conductivity data collected from five Seacat sensors from a mooring as part of the Massachusetts Bay Internal Wave Experiment from 1998-08-05 to 1998-09-01" ;
		:summary = "A 1-month 4-element moored array experiment to measure the currents associated with large-amplitude internal waves generated by tidal flow across Stellwagen Bank" ;
		:source = "WHOI Upper Ocean Proc Grp" ;
		:platform = "mooring, 5391" ;
		:instrument = "Seacat, scat, instrument_1" ;
		:uuid = "" ;
		:sea_name = "Massachusetts Bay, Stellwagen Bank National Marine Sanctuary" ;
		:id = "" ;
		:naming_authority = "gov.noaa.nodc" ;
		:time_coverage_start = "05-Aug-1998 14:46:00" ;
		:time_coverage_end = "01-Sep-1998 16:35:00" ;
		:time_coverage_resolution = "point" ;
		:geospatial_lon_max = -70.3912963867188 ;
		:geospatial_lon_min = -70.3912963867188 ;
		:geospatial_lon_units = "degrees_east" ;
		:geospatial_lon_resolution = "point" ;
		:geospatial_lat_max = 42.3315010070801 ;
		:geospatial_lat_min = 42.3315010070801 ;
		:geospatial_lat_units = "degrees_north" ;
		:geospatial_lat_resolution = "point" ;
		:geospatial_vertical_min = 10. ;
		:geospatial_vertical_max = 50. ;
		:geospatial_vertical_positive = "down" ;
		:geospatial_vertical_units = "meters" ;
		:geospatial_vertical_resolution = "point" ;
		:institution = "U.S.Geological Survey, Woods Hole Coastal and Marine Science Center" ;
		:creator_name = "" ;
		:project = "USGS Coastal Marine Geology Program Sediment Transport group" ;
		:processing_level = "" ;
		:references = "" ;
		:keywords_vocabulary = "" ;
		:keywords = "C:S:T:STH" ;
		:acknowledgment = "original contributor: B. Butman, Project Investigator; data originator: Ellyn Montgomery, WHOI Upper Ocean Proc Grp" ;
		:comment = "" ;
		:contributor_name = "" ;
		:contributor_role = "" ;
		:date_created = "13-Dec-2011" ;
		:date_modified = "13-Dec-2011" ;
		:publisher_name = "US NATIONAL OCEANOGRAPHIC DATA CENTER " ;
		:publisher_email = "NODC.Services@noaa.gov" ;
		:publisher_url = "http://www.nodc.noaa.gov/" ;
		:history = "0 pad values replaced by linear interpolations using EPIC_interp.m :Sample start time fixed.  :Trimmed using truncate.m to select records in the range 3047 to 42036.  :Converted to EPIC by WHOI UOP:, reformatted from EPIC to Climate and Forecast conventions" ;
		:license = "" ;
		:metadata_link = "" ;
}

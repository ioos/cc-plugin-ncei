netcdf wodStandardLevels {
dimensions:
	profile = 169 ;
	z = 26 ;
	strnlen = 170 ;
	strnlensmall = 35 ;
variables:
    int profile(profile) ;
        profile:long_name = "profile long name" ;
        profile:cf_role = "profile_id" ;
	char country(profile, strnlensmall) ;
	char WOD_cruise_identifier(profile, strnlensmall) ;
		WOD_cruise_identifier:comment = "two byte country code + WOD cruise number (unique to country code)" ;
		WOD_cruise_identifier:long_name = "WOD_cruise_identifier" ;
	char originators_cruise_identifier(profile, strnlensmall) ;
	int wod_unique_cast(profile) ;
		wod_unique_cast:cf_role = "profile_id" ;
	char originators_station_identifier(profile, strnlensmall) ;
		originators_station_identifier:long_name = "originators_station_identifier" ;
	float lat(profile) ;
		lat:standard_name = "latitude" ;
		lat:long_name = "latitude" ;
		lat:units = "degrees_north" ;
                lat:axis = "Y" ;
                lat:_FillValue = 0.0f ;
	float lon(profile) ;
		lon:standard_name = "longitude" ;
		lon:long_name = "longitude" ;
		lon:units = "degrees_east" ;
                lon:axis = "X" ;
                lon:_FillValue = 0.0f ;
	double time(profile) ;
		time:standard_name = "time" ;
		time:long_name = "time" ;
		time:units = "days since 1770-01-01 00:00:00" ;
                time:axis = "T" ;
                time:_FillValue = 0.0f ;
                time:calendar = "julian" ;
	int date(profile) ;
		date:long_name = "date" ;
		date:comment = "YYYYMMDD" ;
	float GMT_time(profile) ;
		GMT_time:long_name = "GMT_time" ;
	int Access_no(profile) ;
		Access_no:long_name = "NODC_accession_number" ;
		Access_no:units_wod = "NODC_code" ;
		Access_no:comment = "used to find original data at NODC" ;
	char Project(profile, strnlen) ;
		Project:long_name = "Project_name" ;
		Project:comment = "name or acronym of project under which data were measured" ;
	char Platform(profile, strnlen) ;
		Platform:long_name = "Platform_name" ;
		Platform:comment = "name of platform from which measurements were taken" ;
	char Institute(profile, strnlen) ;
		Institute:long_name = "Responsible_institute" ;
		Institute:comment = "name of institute which collected data" ;
	float Orig_Stat_Num(profile) ;
		Orig_Stat_Num:long_name = "Originators_Station_Number" ;
		Orig_Stat_Num:comment = "number assigned to a given station by data originator" ;
	float Bottom_Depth(profile) ;
		Bottom_Depth:long_name = "Bottom_Depth" ;
		Bottom_Depth:units = "meters" ;
	float Cast_Duration(profile) ;
		Cast_Duration:long_name = "Cast_Duration" ;
		Cast_Duration:units = "hours" ;
	char Water_Color(profile, strnlen) ;
		Water_Color:long_name = "Water_Color" ;
		Water_Color:units_wod = "Forel-Ule scale (00 to 21)" ;
	float Water_Transpar(profile) ;
		Water_Transpar:long_name = "Water_Transparency" ;
		Water_Transpar:units = "meters" ;
		Water_Transpar:comment = "Secchi disk depth" ;
	char Wave_Direction(profile, strnlen) ;
		Wave_Direction:long_name = "Wave_Direction" ;
		Wave_Direction:units_wod = "WMO 0877 or NODC 0110" ;
	char Wave_Height(profile, strnlen) ;
		Wave_Height:long_name = "Wave_Height" ;
		Wave_Height:units_wod = "WMO 1555 or NODC 0104" ;
	char Sea_State(profile, strnlen) ;
		Sea_State:long_name = "Sea_State" ;
		Sea_State:units_wod = "WMO 3700 or NODC 0109" ;
	char Wind_Force(profile, strnlen) ;
		Wind_Force:long_name = "Wind_Force" ;
		Wind_Force:units_wod = "Beaufort scale or NODC 0052" ;
	char Wave_Period(profile, strnlen) ;
		Wave_Period:long_name = "Wave_Period" ;
		Wave_Period:units_wod = "WMO 3155 or NODC 0378" ;
	char Wind_Direction(profile, strnlen) ;
		Wind_Direction:long_name = "Wind_Direction" ;
		Wind_Direction:units_wod = "WMO 0877 or NODC 0110" ;
	float Wind_Speed(profile) ;
		Wind_Speed:long_name = "Wind_Speed" ;
		Wind_Speed:units = "knots" ;
	float Barometric_Pres(profile) ;
		Barometric_Pres:long_name = "Barometric_Pressure" ;
		Barometric_Pres:units = "millibars" ;
	float Dry_Bulb_Temp(profile) ;
		Dry_Bulb_Temp:long_name = "Dry_Bulb_Air_Temperature" ;
		Dry_Bulb_Temp:units = "degree_C" ;
	char Weather_Condition(profile, strnlen) ;
		Weather_Condition:long_name = "Weather_Condition" ;
		Weather_Condition:comment = "Weather conditions at time of measurements" ;
	char Cloud_Type(profile, strnlen) ;
		Cloud_Type:long_name = "Cloud_Type" ;
		Cloud_Type:units_wod = "WMO 0500 or NODC 0053" ;
	char Cloud_Cover(profile, strnlen) ;
		Cloud_Cover:long_name = "Cloud_Cover" ;
		Cloud_Cover:units_wod = "WMO 2700 or NODC 0105" ;
	char dataset(profile, strnlen) ;
		dataset:long_name = "WOD_dataset" ;
	char Ref_Type(profile, strnlen) ;
		Ref_Type:long_name = "Reference_Instrument" ;
		Ref_Type:comment = "Instrument for reference temperature" ;
	char Visibility(profile, strnlen) ;
		Visibility:long_name = "Horizontal_visibility" ;
		Visibility:units_wod = "WMO Code 4300" ;
	float Absol_Humidity(profile) ;
		Absol_Humidity:long_name = "Absolute_Humidity" ;
		Absol_Humidity:units = "gram/m3" ;
	char dbase_orig(profile, strnlen) ;
		dbase_orig:long_name = "database_origin" ;
		dbase_orig:comment = "Database from which data were extracted" ;
	float z(z) ;
		z:standard_name = "altitude" ;
		z:long_name = "depth_below_sea_level" ;
		z:units = "m" ;
		z:positive = "down" ;
                z:axis = "Z" ;
	short zcast_WODflag(profile, z) ;
		zcast_WODflag:flag_definitions = "WODfd" ;
	float Temperature(profile, z) ;
		Temperature:long_name = "Temperature" ;
		Temperature:standard_name = "sea_water_temperature" ;
		Temperature:units = "degree_C" ;
		Temperature:coordinates = "time lat lon z" ;
		Temperature:grid_mapping = "crs" ;
	short Temperature_sigfigs(profile, z) ;
	short Temperature_WODflag(profile, z) ;
		Temperature_WODflag:flag_definitions = "WODf" ;
	short Temperature_WODprofileflag(profile) ;
		Temperature_WODprofileflag:flag_definitions = "WODfp" ;
	char Temperature_Instrument(profile, strnlen) ;
		Temperature_Instrument:long_name = "Instrument" ;
		Temperature_Instrument:comment = "Device used for measurement" ;
	float Salinity(profile, z) ;
		Salinity:long_name = "Salinity" ;
		Salinity:standard_name = "sea_water_salinity" ;
		Salinity:coordinates = "time lat lon z" ;
		Salinity:grid_mapping = "crs" ;
	short Salinity_sigfigs(profile, z) ;
	short Salinity_WODflag(profile, z) ;
		Salinity_WODflag:flag_definitions = "WODf" ;
	short Salinity_WODprofileflag(profile) ;
		Salinity_WODprofileflag:flag_definitions = "WODfp" ;
	char Salinity_Instrument(profile, strnlen) ;
		Salinity_Instrument:long_name = "Instrument" ;
		Salinity_Instrument:comment = "Device used for measurement" ;
	float Oxygen(profile, z) ;
		Oxygen:long_name = "Oxygen" ;
		Oxygen:standard_name = "volume_fraction_of_oxygen_in_sea_water" ;
		Oxygen:units = "ml/l" ;
		Oxygen:coordinates = "time lat lon z" ;
		Oxygen:grid_mapping = "crs" ;
	short Oxygen_sigfigs(profile, z) ;
	short Oxygen_WODflag(profile, z) ;
		Oxygen_WODflag:flag_definitions = "WODf" ;
	short Oxygen_WODprofileflag(profile) ;
		Oxygen_WODprofileflag:flag_definitions = "WODfp" ;
	char Oxygen_Original_units(profile, strnlen) ;
		Oxygen_Original_units:comment = "Units originally used: coverted to standard units" ;
	float Phosphate(profile, z) ;
		Phosphate:long_name = "Phosphate" ;
		Phosphate:standard_name = "mole_concentration_of_phosphate_in_sea_water" ;
		Phosphate:units = "umol/l" ;
		Phosphate:coordinates = "time lat lon z" ;
		Phosphate:grid_mapping = "crs" ;
	short Phosphate_sigfigs(profile, z) ;
	short Phosphate_WODflag(profile, z) ;
		Phosphate_WODflag:flag_definitions = "WODf" ;
	short Phosphate_WODprofileflag(profile) ;
		Phosphate_WODprofileflag:flag_definitions = "WODfp" ;
	char Phosphate_Original_units(profile, strnlen) ;
		Phosphate_Original_units:comment = "Units originally used: coverted to standard units" ;
	float TotalPhos(profile, z) ;
		TotalPhos:long_name = "TotalPhos" ;
		TotalPhos:units = "umol/l" ;
		TotalPhos:coordinates = "time lat lon z" ;
		TotalPhos:grid_mapping = "crs" ;
	short TotalPhos_sigfigs(profile, z) ;
	short TotalPhos_WODflag(profile, z) ;
		TotalPhos_WODflag:flag_definitions = "WODf" ;
	float Silicate(profile, z) ;
		Silicate:long_name = "Silicate" ;
		Silicate:standard_name = "mole_concentration_of_silicate_in_sea_water" ;
		Silicate:units = "umol/l" ;
		Silicate:coordinates = "time lat lon z" ;
		Silicate:grid_mapping = "crs" ;
	short Silicate_sigfigs(profile, z) ;
	short Silicate_WODflag(profile, z) ;
		Silicate_WODflag:flag_definitions = "WODf" ;
	short Silicate_WODprofileflag(profile) ;
		Silicate_WODprofileflag:flag_definitions = "WODfp" ;
	char Silicate_Original_units(profile, strnlen) ;
		Silicate_Original_units:comment = "Units originally used: coverted to standard units" ;
	float Nitrite(profile, z) ;
		Nitrite:long_name = "Nitrite" ;
		Nitrite:units = "umol/l" ;
		Nitrite:coordinates = "time lat lon z" ;
		Nitrite:grid_mapping = "crs" ;
	short Nitrite_sigfigs(profile, z) ;
	short Nitrite_WODflag(profile, z) ;
		Nitrite_WODflag:flag_definitions = "WODf" ;
	char Nitrite_Original_units(profile, strnlen) ;
		Nitrite_Original_units:comment = "Units originally used: coverted to standard units" ;
	float Nitrate(profile, z) ;
		Nitrate:long_name = "Nitrate" ;
		Nitrate:standard_name = "mole_concentration_of_nitrate_in_sea_water" ;
		Nitrate:units = "umol/l" ;
		Nitrate:coordinates = "time lat lon z" ;
		Nitrate:grid_mapping = "crs" ;
	short Nitrate_sigfigs(profile, z) ;
	short Nitrate_WODflag(profile, z) ;
		Nitrate_WODflag:flag_definitions = "WODf" ;
	short Nitrate_WODprofileflag(profile) ;
		Nitrate_WODprofileflag:flag_definitions = "WODfp" ;
	char Nitrate_Original_units(profile, strnlen) ;
		Nitrate_Original_units:comment = "Units originally used: coverted to standard units" ;
	float pH(profile, z) ;
		pH:long_name = "sea_water_ph" ;
		pH:coordinates = "time lat lon z" ;
		pH:grid_mapping = "crs" ;
	short pH_sigfigs(profile, z) ;
	short pH_WODflag(profile, z) ;
		pH_WODflag:flag_definitions = "WODf" ;
	short pH_WODprofileflag(profile) ;
		pH_WODprofileflag:flag_definitions = "WODfp" ;
	float Ammonia(profile, z) ;
		Ammonia:long_name = "Ammonia" ;
		Ammonia:coordinates = "time lat lon z" ;
		Ammonia:grid_mapping = "crs" ;
	short Ammonia_sigfigs(profile, z) ;
	short Ammonia_WODflag(profile, z) ;
		Ammonia_WODflag:flag_definitions = "WODf" ;
	float Chlorophyll(profile, z) ;
		Chlorophyll:long_name = "Chlorophyll" ;
		Chlorophyll:standard_name = "mass_concentration_of_chlorophyll_in_sea_water" ;
		Chlorophyll:units = "ugram/l" ;
		Chlorophyll:coordinates = "time lat lon z" ;
		Chlorophyll:grid_mapping = "crs" ;
	short Chlorophyll_sigfigs(profile, z) ;
	short Chlorophyll_WODflag(profile, z) ;
		Chlorophyll_WODflag:flag_definitions = "WODf" ;
	short Chlorophyll_WODprofileflag(profile) ;
		Chlorophyll_WODprofileflag:flag_definitions = "WODfp" ;
	float Phaeophytin(profile, z) ;
		Phaeophytin:long_name = "Phaeophytin" ;
		Phaeophytin:coordinates = "time lat lon z" ;
		Phaeophytin:grid_mapping = "crs" ;
	short Phaeophytin_sigfigs(profile, z) ;
	short Phaeophytin_WODflag(profile, z) ;
		Phaeophytin_WODflag:flag_definitions = "WODf" ;
	float Alkalinity(profile, z) ;
		Alkalinity:long_name = "Alkalinity" ;
		Alkalinity:standard_name = "sea_water_alkalinity_expressed_as_mole_equivalent" ;
		Alkalinity:units = "umol/l" ;
		Alkalinity:coordinates = "time lat lon z" ;
		Alkalinity:grid_mapping = "crs" ;
	short Alkalinity_sigfigs(profile, z) ;
	short Alkalinity_WODflag(profile, z) ;
		Alkalinity_WODflag:flag_definitions = "WODf" ;
	short Alkalinity_WODprofileflag(profile) ;
		Alkalinity_WODprofileflag:flag_definitions = "WODfp" ;
	float NO2NO3(profile, z) ;
		NO2NO3:long_name = "NO2NO3" ;
		NO2NO3:units = "umol/l" ;
		NO2NO3:coordinates = "time lat lon z" ;
		NO2NO3:grid_mapping = "crs" ;
	short NO2NO3_sigfigs(profile, z) ;
	short NO2NO3_WODflag(profile, z) ;
		NO2NO3_WODflag:flag_definitions = "WODf" ;
	int crs ;
		crs:grid_mapping_name = "latitude_longitude" ;
		crs:epsg_code = "EPSG:4326" ;
		crs:longitude_of_prime_meridian = 0.f ;
		crs:semi_major_axis = 6378137.f ;
		crs:inverse_flattening = 298.2572f ;
	short WODf ;
		WODf:long_name = "WOD_standard_level_flag" ;
		WODf:flag_values = 0s, 1s, 2s, 3s, 4s, 5s, 6s, 7s, 8s, 9s ;
		WODf:flag_meanings = "accepted anomaly density_inversion annual_sd_out seasonal_sd_out monthly_sd_out annual+seasonal_sd_out annual+monthly_sd_out seasonal+monthly_sd_out annual+seasonal+monthly_sd_out" ;
	short WODfp ;
		WODfp:long_name = "WOD_profile_flag" ;
		WODfp:flag_values = 0s, 1s, 2s, 3s, 4s, 5s, 6s, 7s, 8s, 9s ;
		WODfp:flag_meanings = "accepted annual_sd_out density_inversion cruise seasonal_sd_out monthly_sd_out annual+seasonal_sd_out anomaly_or_annual+monthly_sd_out seasonal+monthly_sd_out annual+seasonal+monthly_sd_out" ;
	short WODfd ;
		WODfd:long_name = "WOD_depth_level_" ;
		WODfd:flag_values = 0s, 1s, 2s ;
		WODfd:flag_meanings = "accepted duplicate_or_inversion density_inversion" ;

// global attributes:
		:standard_name_vocabulary = "NetCDF Climate and Forecast (CF) Metadata Convention Standard Name Table v23" ;
		:featureType = "profile" ;
		:cdm_data_type = "Station" ;
		:Conventions = "CF-1.6" ;
                :Metadata_Conventions = "Unidata Dataset Discovery v1.0" ;
                :nodc_template_version = "NODC_NetCDF_Profile_Orthogonal_Template_v1.1" ;
}

netcdf wodStandardLevels {
dimensions:
	profile = 169 ;
	z = 26 ;
	strnlen = 170 ;
	strnlensmall = 35 ;
variables:
    int profile(profile) ;
        profile:long_name = "profile long name" ;
        profile:cf_role = "profile_id" ;
	char country(profile, strnlensmall) ;
	char WOD_cruise_identifier(profile, strnlensmall) ;
		WOD_cruise_identifier:comment = "two byte country code + WOD cruise number (unique to country code)" ;
		WOD_cruise_identifier:long_name = "WOD_cruise_identifier" ;
	char originators_cruise_identifier(profile, strnlensmall) ;
	int wod_unique_cast(profile) ;
		wod_unique_cast:cf_role = "profile_id" ;
	char originators_station_identifier(profile, strnlensmall) ;
		originators_station_identifier:long_name = "originators_station_identifier" ;
	float lat(profile) ;
		lat:standard_name = "latitude" ;
		lat:long_name = "latitude" ;
		lat:units = "degrees_north" ;
                lat:axis = "Y" ;
                lat:_FillValue = 0.0f ;
	float lon(profile) ;
		lon:standard_name = "longitude" ;
		lon:long_name = "longitude" ;
		lon:units = "degrees_east" ;
                lon:axis = "X" ;
                lon:_FillValue = 0.0f ;
	double time(profile) ;
		time:standard_name = "time" ;
		time:long_name = "time" ;
		time:units = "days since 1770-01-01 00:00:00" ;
                time:axis = "T" ;
                time:_FillValue = 0.0f ;
                time:calendar = "julian" ;
	int date(profile) ;
		date:long_name = "date" ;
		date:comment = "YYYYMMDD" ;
	float GMT_time(profile) ;
		GMT_time:long_name = "GMT_time" ;
	int Access_no(profile) ;
		Access_no:long_name = "NODC_accession_number" ;
		Access_no:units_wod = "NODC_code" ;
		Access_no:comment = "used to find original data at NODC" ;
	char Project(profile, strnlen) ;
		Project:long_name = "Project_name" ;
		Project:comment = "name or acronym of project under which data were measured" ;
	char Platform(profile, strnlen) ;
		Platform:long_name = "Platform_name" ;
		Platform:comment = "name of platform from which measurements were taken" ;
	char Institute(profile, strnlen) ;
		Institute:long_name = "Responsible_institute" ;
		Institute:comment = "name of institute which collected data" ;
	float Orig_Stat_Num(profile) ;
		Orig_Stat_Num:long_name = "Originators_Station_Number" ;
		Orig_Stat_Num:comment = "number assigned to a given station by data originator" ;
	float Bottom_Depth(profile) ;
		Bottom_Depth:long_name = "Bottom_Depth" ;
		Bottom_Depth:units = "meters" ;
	float Cast_Duration(profile) ;
		Cast_Duration:long_name = "Cast_Duration" ;
		Cast_Duration:units = "hours" ;
	char Water_Color(profile, strnlen) ;
		Water_Color:long_name = "Water_Color" ;
		Water_Color:units_wod = "Forel-Ule scale (00 to 21)" ;
	float Water_Transpar(profile) ;
		Water_Transpar:long_name = "Water_Transparency" ;
		Water_Transpar:units = "meters" ;
		Water_Transpar:comment = "Secchi disk depth" ;
	char Wave_Direction(profile, strnlen) ;
		Wave_Direction:long_name = "Wave_Direction" ;
		Wave_Direction:units_wod = "WMO 0877 or NODC 0110" ;
	char Wave_Height(profile, strnlen) ;
		Wave_Height:long_name = "Wave_Height" ;
		Wave_Height:units_wod = "WMO 1555 or NODC 0104" ;
	char Sea_State(profile, strnlen) ;
		Sea_State:long_name = "Sea_State" ;
		Sea_State:units_wod = "WMO 3700 or NODC 0109" ;
	char Wind_Force(profile, strnlen) ;
		Wind_Force:long_name = "Wind_Force" ;
		Wind_Force:units_wod = "Beaufort scale or NODC 0052" ;
	char Wave_Period(profile, strnlen) ;
		Wave_Period:long_name = "Wave_Period" ;
		Wave_Period:units_wod = "WMO 3155 or NODC 0378" ;
	char Wind_Direction(profile, strnlen) ;
		Wind_Direction:long_name = "Wind_Direction" ;
		Wind_Direction:units_wod = "WMO 0877 or NODC 0110" ;
	float Wind_Speed(profile) ;
		Wind_Speed:long_name = "Wind_Speed" ;
		Wind_Speed:units = "knots" ;
	float Barometric_Pres(profile) ;
		Barometric_Pres:long_name = "Barometric_Pressure" ;
		Barometric_Pres:units = "millibars" ;
	float Dry_Bulb_Temp(profile) ;
		Dry_Bulb_Temp:long_name = "Dry_Bulb_Air_Temperature" ;
		Dry_Bulb_Temp:units = "degree_C" ;
	char Weather_Condition(profile, strnlen) ;
		Weather_Condition:long_name = "Weather_Condition" ;
		Weather_Condition:comment = "Weather conditions at time of measurements" ;
	char Cloud_Type(profile, strnlen) ;
		Cloud_Type:long_name = "Cloud_Type" ;
		Cloud_Type:units_wod = "WMO 0500 or NODC 0053" ;
	char Cloud_Cover(profile, strnlen) ;
		Cloud_Cover:long_name = "Cloud_Cover" ;
		Cloud_Cover:units_wod = "WMO 2700 or NODC 0105" ;
	char dataset(profile, strnlen) ;
		dataset:long_name = "WOD_dataset" ;
	char Ref_Type(profile, strnlen) ;
		Ref_Type:long_name = "Reference_Instrument" ;
		Ref_Type:comment = "Instrument for reference temperature" ;
	char Visibility(profile, strnlen) ;
		Visibility:long_name = "Horizontal_visibility" ;
		Visibility:units_wod = "WMO Code 4300" ;
	float Absol_Humidity(profile) ;
		Absol_Humidity:long_name = "Absolute_Humidity" ;
		Absol_Humidity:units = "gram/m3" ;
	char dbase_orig(profile, strnlen) ;
		dbase_orig:long_name = "database_origin" ;
		dbase_orig:comment = "Database from which data were extracted" ;
	float z(z) ;
		z:standard_name = "altitude" ;
		z:long_name = "depth_below_sea_level" ;
		z:units = "m" ;
		z:positive = "down" ;
                z:axis = "Z" ;
	short zcast_WODflag(profile, z) ;
		zcast_WODflag:flag_definitions = "WODfd" ;
	float Temperature(profile, z) ;
		Temperature:long_name = "Temperature" ;
		Temperature:standard_name = "sea_water_temperature" ;
		Temperature:units = "degree_C" ;
		Temperature:coordinates = "time lat lon z" ;
		Temperature:grid_mapping = "crs" ;
	short Temperature_sigfigs(profile, z) ;
	short Temperature_WODflag(profile, z) ;
		Temperature_WODflag:flag_definitions = "WODf" ;
	short Temperature_WODprofileflag(profile) ;
		Temperature_WODprofileflag:flag_definitions = "WODfp" ;
	char Temperature_Instrument(profile, strnlen) ;
		Temperature_Instrument:long_name = "Instrument" ;
		Temperature_Instrument:comment = "Device used for measurement" ;
	float Salinity(profile, z) ;
		Salinity:long_name = "Salinity" ;
		Salinity:standard_name = "sea_water_salinity" ;
		Salinity:coordinates = "time lat lon z" ;
		Salinity:grid_mapping = "crs" ;
	short Salinity_sigfigs(profile, z) ;
	short Salinity_WODflag(profile, z) ;
		Salinity_WODflag:flag_definitions = "WODf" ;
	short Salinity_WODprofileflag(profile) ;
		Salinity_WODprofileflag:flag_definitions = "WODfp" ;
	char Salinity_Instrument(profile, strnlen) ;
		Salinity_Instrument:long_name = "Instrument" ;
		Salinity_Instrument:comment = "Device used for measurement" ;
	float Oxygen(profile, z) ;
		Oxygen:long_name = "Oxygen" ;
		Oxygen:standard_name = "volume_fraction_of_oxygen_in_sea_water" ;
		Oxygen:units = "ml/l" ;
		Oxygen:coordinates = "time lat lon z" ;
		Oxygen:grid_mapping = "crs" ;
	short Oxygen_sigfigs(profile, z) ;
	short Oxygen_WODflag(profile, z) ;
		Oxygen_WODflag:flag_definitions = "WODf" ;
	short Oxygen_WODprofileflag(profile) ;
		Oxygen_WODprofileflag:flag_definitions = "WODfp" ;
	char Oxygen_Original_units(profile, strnlen) ;
		Oxygen_Original_units:comment = "Units originally used: coverted to standard units" ;
	float Phosphate(profile, z) ;
		Phosphate:long_name = "Phosphate" ;
		Phosphate:standard_name = "mole_concentration_of_phosphate_in_sea_water" ;
		Phosphate:units = "umol/l" ;
		Phosphate:coordinates = "time lat lon z" ;
		Phosphate:grid_mapping = "crs" ;
	short Phosphate_sigfigs(profile, z) ;
	short Phosphate_WODflag(profile, z) ;
		Phosphate_WODflag:flag_definitions = "WODf" ;
	short Phosphate_WODprofileflag(profile) ;
		Phosphate_WODprofileflag:flag_definitions = "WODfp" ;
	char Phosphate_Original_units(profile, strnlen) ;
		Phosphate_Original_units:comment = "Units originally used: coverted to standard units" ;
	float TotalPhos(profile, z) ;
		TotalPhos:long_name = "TotalPhos" ;
		TotalPhos:units = "umol/l" ;
		TotalPhos:coordinates = "time lat lon z" ;
		TotalPhos:grid_mapping = "crs" ;
	short TotalPhos_sigfigs(profile, z) ;
	short TotalPhos_WODflag(profile, z) ;
		TotalPhos_WODflag:flag_definitions = "WODf" ;
	float Silicate(profile, z) ;
		Silicate:long_name = "Silicate" ;
		Silicate:standard_name = "mole_concentration_of_silicate_in_sea_water" ;
		Silicate:units = "umol/l" ;
		Silicate:coordinates = "time lat lon z" ;
		Silicate:grid_mapping = "crs" ;
	short Silicate_sigfigs(profile, z) ;
	short Silicate_WODflag(profile, z) ;
		Silicate_WODflag:flag_definitions = "WODf" ;
	short Silicate_WODprofileflag(profile) ;
		Silicate_WODprofileflag:flag_definitions = "WODfp" ;
	char Silicate_Original_units(profile, strnlen) ;
		Silicate_Original_units:comment = "Units originally used: coverted to standard units" ;
	float Nitrite(profile, z) ;
		Nitrite:long_name = "Nitrite" ;
		Nitrite:units = "umol/l" ;
		Nitrite:coordinates = "time lat lon z" ;
		Nitrite:grid_mapping = "crs" ;
	short Nitrite_sigfigs(profile, z) ;
	short Nitrite_WODflag(profile, z) ;
		Nitrite_WODflag:flag_definitions = "WODf" ;
	char Nitrite_Original_units(profile, strnlen) ;
		Nitrite_Original_units:comment = "Units originally used: coverted to standard units" ;
	float Nitrate(profile, z) ;
		Nitrate:long_name = "Nitrate" ;
		Nitrate:standard_name = "mole_concentration_of_nitrate_in_sea_water" ;
		Nitrate:units = "umol/l" ;
		Nitrate:coordinates = "time lat lon z" ;
		Nitrate:grid_mapping = "crs" ;
	short Nitrate_sigfigs(profile, z) ;
	short Nitrate_WODflag(profile, z) ;
		Nitrate_WODflag:flag_definitions = "WODf" ;
	short Nitrate_WODprofileflag(profile) ;
		Nitrate_WODprofileflag:flag_definitions = "WODfp" ;
	char Nitrate_Original_units(profile, strnlen) ;
		Nitrate_Original_units:comment = "Units originally used: coverted to standard units" ;
	float pH(profile, z) ;
		pH:long_name = "sea_water_ph" ;
		pH:coordinates = "time lat lon z" ;
		pH:grid_mapping = "crs" ;
	short pH_sigfigs(profile, z) ;
	short pH_WODflag(profile, z) ;
		pH_WODflag:flag_definitions = "WODf" ;
	short pH_WODprofileflag(profile) ;
		pH_WODprofileflag:flag_definitions = "WODfp" ;
	float Ammonia(profile, z) ;
		Ammonia:long_name = "Ammonia" ;
		Ammonia:coordinates = "time lat lon z" ;
		Ammonia:grid_mapping = "crs" ;
	short Ammonia_sigfigs(profile, z) ;
	short Ammonia_WODflag(profile, z) ;
		Ammonia_WODflag:flag_definitions = "WODf" ;
	float Chlorophyll(profile, z) ;
		Chlorophyll:long_name = "Chlorophyll" ;
		Chlorophyll:standard_name = "mass_concentration_of_chlorophyll_in_sea_water" ;
		Chlorophyll:units = "ugram/l" ;
		Chlorophyll:coordinates = "time lat lon z" ;
		Chlorophyll:grid_mapping = "crs" ;
	short Chlorophyll_sigfigs(profile, z) ;
	short Chlorophyll_WODflag(profile, z) ;
		Chlorophyll_WODflag:flag_definitions = "WODf" ;
	short Chlorophyll_WODprofileflag(profile) ;
		Chlorophyll_WODprofileflag:flag_definitions = "WODfp" ;
	float Phaeophytin(profile, z) ;
		Phaeophytin:long_name = "Phaeophytin" ;
		Phaeophytin:coordinates = "time lat lon z" ;
		Phaeophytin:grid_mapping = "crs" ;
	short Phaeophytin_sigfigs(profile, z) ;
	short Phaeophytin_WODflag(profile, z) ;
		Phaeophytin_WODflag:flag_definitions = "WODf" ;
	float Alkalinity(profile, z) ;
		Alkalinity:long_name = "Alkalinity" ;
		Alkalinity:standard_name = "sea_water_alkalinity_expressed_as_mole_equivalent" ;
		Alkalinity:units = "umol/l" ;
		Alkalinity:coordinates = "time lat lon z" ;
		Alkalinity:grid_mapping = "crs" ;
	short Alkalinity_sigfigs(profile, z) ;
	short Alkalinity_WODflag(profile, z) ;
		Alkalinity_WODflag:flag_definitions = "WODf" ;
	short Alkalinity_WODprofileflag(profile) ;
		Alkalinity_WODprofileflag:flag_definitions = "WODfp" ;
	float NO2NO3(profile, z) ;
		NO2NO3:long_name = "NO2NO3" ;
		NO2NO3:units = "umol/l" ;
		NO2NO3:coordinates = "time lat lon z" ;
		NO2NO3:grid_mapping = "crs" ;
	short NO2NO3_sigfigs(profile, z) ;
	short NO2NO3_WODflag(profile, z) ;
		NO2NO3_WODflag:flag_definitions = "WODf" ;
	int crs ;
		crs:grid_mapping_name = "latitude_longitude" ;
		crs:epsg_code = "EPSG:4326" ;
		crs:longitude_of_prime_meridian = 0.f ;
		crs:semi_major_axis = 6378137.f ;
		crs:inverse_flattening = 298.2572f ;
	short WODf ;
		WODf:long_name = "WOD_standard_level_flag" ;
		WODf:flag_values = 0s, 1s, 2s, 3s, 4s, 5s, 6s, 7s, 8s, 9s ;
		WODf:flag_meanings = "accepted anomaly density_inversion annual_sd_out seasonal_sd_out monthly_sd_out annual+seasonal_sd_out annual+monthly_sd_out seasonal+monthly_sd_out annual+seasonal+monthly_sd_out" ;
	short WODfp ;
		WODfp:long_name = "WOD_profile_flag" ;
		WODfp:flag_values = 0s, 1s, 2s, 3s, 4s, 5s, 6s, 7s, 8s, 9s ;
		WODfp:flag_meanings = "accepted annual_sd_out density_inversion cruise seasonal_sd_out monthly_sd_out annual+seasonal_sd_out anomaly_or_annual+monthly_sd_out seasonal+monthly_sd_out annual+seasonal+monthly_sd_out" ;
	short WODfd ;
		WODfd:long_name = "WOD_depth_level_" ;
		WODfd:flag_values = 0s, 1s, 2s ;
		WODfd:flag_meanings = "accepted duplicate_or_inversion density_inversion" ;

// global attributes:
		:standard_name_vocabulary = "NetCDF Climate and Forecast (CF) Metadata Convention Standard Name Table v23" ;
		:featureType = "profile" ;
		:cdm_data_type = "Station" ;
		:Conventions = "CF-1.6" ;
                :Metadata_Conventions = "Unidata Dataset Discovery v1.0" ;
                :nodc_template_version = "NODC_NetCDF_Profile_Orthogonal_Template_v1.1" ;
data:

 country =
  "JAPAN",
  "SOVIET UNION",
  "CANADA",
  "UNITED STATES",
  "POLAND",
  "SOVIET UNION",
  "NORWAY",
  "JAPAN",
  "CANADA",
  "CANADA",
  "NORWAY",
  "SOVIET UNION",
  "CANADA",
  "NORWAY",
  "JAPAN",
  "SOVIET UNION",
  "SOVIET UNION",
  "CANADA",
  "UNITED STATES",
  "SOVIET UNION",
  "JAPAN",
  "NORWAY",
  "CANADA",
  "UNITED STATES",
  "SOVIET UNION",
  "SOVIET UNION",
  "CANADA",
  "NORWAY",
  "SOVIET UNION",
  "NORWAY",
  "POLAND",
  "JAPAN",
  "JAPAN",
  "UNITED STATES",
  "NORWAY",
  "JAPAN",
  "SOVIET UNION",
  "SOVIET UNION",
  "CANADA",
  "JAPAN",
  "SOVIET UNION",
  "NORWAY",
  "CANADA",
  "SOVIET UNION",
  "GREAT BRITAIN",
  "GREAT BRITAIN",
  "NORWAY",
  "CANADA",
  "SOVIET UNION",
  "SOVIET UNION",
  "SOVIET UNION",
  "GREAT BRITAIN",
  "POLAND",
  "UNITED STATES",
  "NORWAY",
  "CANADA",
  "UNITED STATES",
  "NORWAY",
  "SOVIET UNION",
  "NORWAY",
  "UNITED STATES",
  "GREAT BRITAIN",
  "GREAT BRITAIN",
  "SOVIET UNION",
  "NETHERLANDS",
  "NORWAY",
  "CANADA",
  "CANADA",
  "FRANCE",
  "SOVIET UNION",
  "GREAT BRITAIN",
  "BELGIUM",
  "NORWAY",
  "GREAT BRITAIN",
  "CANADA",
  "SOVIET UNION",
  "CANADA",
  "POLAND",
  "UNITED STATES",
  "EAST GERMANY",
  "NORWAY",
  "UNITED STATES",
  "UNITED STATES",
  "GREAT BRITAIN",
  "JAPAN",
  "NORWAY",
  "SOVIET UNION",
  "SOVIET UNION",
  "SOVIET UNION",
  "CANADA",
  "SOVIET UNION",
  "SOVIET UNION",
  "NORWAY",
  "BELGIUM",
  "CANADA",
  "SOVIET UNION",
  "SOVIET UNION",
  "SOVIET UNION",
  "SOVIET UNION",
  "NORWAY",
  "NORWAY",
  "BELGIUM",
  "SOVIET UNION",
  "SOVIET UNION",
  "NORWAY",
  "NORWAY",
  "BELGIUM",
  "SOVIET UNION",
  "EAST GERMANY",
  "CANADA",
  "UNITED STATES",
  "SOVIET UNION",
  "POLAND",
  "SOVIET UNION",
  "NORWAY",
  "CANADA",
  "BELGIUM",
  "UNITED STATES",
  "EAST GERMANY",
  "NORWAY",
  "NORWAY",
  "CANADA",
  "JAPAN",
  "UNITED STATES",
  "SOVIET UNION",
  "SOVIET UNION",
  "SOVIET UNION",
  "CANADA",
  "UNITED STATES",
  "UNITED STATES",
  "NORWAY",
  "BELGIUM",
  "BELGIUM",
  "UNITED STATES",
  "CANADA",
  "SOVIET UNION",
  "EAST GERMANY",
  "NORWAY",
  "SOVIET UNION",
  "SOVIET UNION",
  "SOVIET UNION",
  "CANADA",
  "UNITED STATES",
  "CANADA",
  "EAST GERMANY",
  "CANADA",
  "UNITED STATES",
  "SOVIET UNION",
  "CANADA",
  "CANADA",
  "UNITED STATES",
  "JAPAN",
  "CANADA",
  "SOVIET UNION",
  "SOVIET UNION",
  "UNITED STATES",
  "NORWAY",
  "SOVIET UNION",
  "GREAT BRITAIN",
  "GREAT BRITAIN",
  "AUSTRALIA",
  "GREAT BRITAIN",
  "UNITED STATES",
  "GREAT BRITAIN",
  "CANADA",
  "GREAT BRITAIN",
  "GREAT BRITAIN",
  "GREAT BRITAIN",
  "GREAT BRITAIN" ;

 WOD_cruise_identifier =
  "JP014480",
  "SU000710",
  "CA001266",
  "US003039",
  "PL000108",
  "SU007601",
  "NO001925",
  "JP026717",
  "CA001267",
  "CA012236",
  "NO001924",
  "SU015381",
  "CA001266",
  "NO001925",
  "JP026717",
  "SU000712",
  "SU015255",
  "CA001266",
  "US003039",
  "SU000713",
  "JP026717",
  "NO001924",
  "CA001267",
  "US003039",
  "SU015463",
  "SU017947",
  "CA001266",
  "NO001925",
  "SU008680",
  "NO001925",
  "PL000108",
  "JP026717",
  "JP026717",
  "US010256",
  "NO001925",
  "JP026717",
  "SU015256",
  "SU017948",
  "CA001266",
  "JP014480",
  "SU000710",
  "NO001132",
  "CA001267",
  "SU007601",
  "GB009271",
  "GB009271",
  "NO001132",
  "CA001266",
  "SU000712",
  "SU017947",
  "SU015255",
  "GB009271",
  "PL000108",
  "US003039",
  "NO001925",
  "CA001266",
  "US003039",
  "NO001924",
  "SU008680",
  "NO001926",
  "US010256",
  "GB009271",
  "GB009271",
  "SU015463",
  "NL001252",
  "NO001926",
  "CA001267",
  "CA001266",
  "FR008171",
  "SU014053",
  "GB009271",
  "BE001100",
  "NO001926",
  "GB009271",
  "CA001266",
  "SU015256",
  "CA001267",
  "PL000108",
  "US003039",
  "DU000339",
  "NO001925",
  "US003039",
  "US010256",
  "GB009271",
  "JP014480",
  "NO001926",
  "SU008678",
  "SU017948",
  "SU015255",
  "CA001267",
  "SU000722",
  "SU007825",
  "NO001925",
  "BE001100",
  "CA001266",
  "SU015463",
  "SU007601",
  "SU021561",
  "SU021561",
  "NO001924",
  "NO001926",
  "BE001100",
  "SU008680",
  "SU021561",
  "NO001925",
  "NO001924",
  "BE001100",
  "SU000712",
  "DU000339",
  "CA001266",
  "US010256",
  "SU000713",
  "PL000108",
  "SU015256",
  "NO001926",
  "CA001266",
  "BE001100",
  "US003039",
  "DU000339",
  "NO001924",
  "NO001926",
  "CA001267",
  "JP014480",
  "US003039",
  "SU007825",
  "SU015463",
  "SU015255",
  "CA001266",
  "US003039",
  "US003039",
  "NO001926",
  "BE001100",
  "BE001100",
  "US008606",
  "CA001267",
  "SU008680",
  "DU000339",
  "NO001926",
  "SU015256",
  "SU007601",
  "SU015255",
  "CA001266",
  "US003039",
  "CA001267",
  "DU000339",
  "CA001266",
  "US003039",
  "SU015463",
  "CA001266",
  "CA001266",
  "US003039",
  "JP014480",
  "CA001267",
  "SU007091",
  "SU015255",
  "US003039",
  "NO001924",
  "SU008680",
  "GB009270",
  "GB009270",
  "AU002470",
  "GB009270",
  "US010724",
  "GB009270",
  "CA008597",
  "GB009270",
  "GB009270",
  "GB009270",
  "GB009270" ;

 originators_cruise_identifier =
  "26",
  "18038000",
  "AL8002",
  "80-02",
  "4",
  "_US2_1980 06",
  "18038000",
  "80003",
  "8",
  "18038000",
  "_US2_1980 06",
  "25",
  "9",
  "18038000",
  "AL8002",
  "33",
  "_US2_1980 06",
  "18038000",
  "AL8002",
  "28",
  "18038000",
  "25",
  "80-02",
  "_US2_1980 06",
  "_US2_1980 06",
  "WI8002",
  "_US2_1980 06",
  "18038000",
  "26",
  "18038000",
  "4",
  "18038000",
  "25",
  "9",
  "80-02",
  "AL8002",
  "18038000",
  "AL8002",
  "25",
  "WI8002",
  "28",
  "18038000",
  "18038000",
  "BN809000",
  "3",
  "18038000",
  "18038000",
  "80-02",
  "AL8002",
  "AL8002",
  "WI8002",
  "19",
  "9",
  "18038000",
  "31",
  "18038000",
  "28",
  "4",
  "25",
  "25",
  "18038000",
  "WI8002",
  "33",
  "80-02",
  "18038000",
  "AL8002",
  "18038000",
  "AL8002",
  "28",
  "9",
  "18038000",
  "AL8002",
  "AL8002",
  "002",
  "18038000",
  "25",
  "4",
  "9",
  "18038000",
  "AL8002",
  "18038000",
  "18038000",
  "AL8002",
  "28",
  "18038000",
  "18038000",
  "AL8002",
  "18038000",
  "26",
  "9",
  "AL8002",
  "25",
  "OWS PAPA",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "" ;

 wod_unique_cast = 7939893, 788994, 788996, 788995, 11119672, 10253223, 
    6876518, 8933719, 788998, 6876515, 6876517, 9966443, 788999, 6876519, 
    8933720, 789000, 9640274, 789002, 6876468, 789003, 8933721, 6876521, 
    789004, 789001, 9977033, 11239237, 789006, 6876524, 6876525, 6876526, 
    789005, 8933723, 8933722, 6876474, 6876527, 8933724, 9966444, 11239238, 
    789007, 7939894, 789009, 6876529, 789008, 10253224, 6876533, 6876534, 
    6876535, 789010, 789011, 11239239, 9640275, 6876542, 789014, 789012, 
    6876537, 789013, 6876481, 6876540, 6876536, 6876538, 6876483, 6876539, 
    6876541, 9977034, 6876543, 6876545, 789016, 789015, 789018, 8553281, 
    6876547, 7732815, 6876548, 6876550, 789017, 9966445, 789020, 789021, 
    789019, 6876557, 6876555, 7506022, 6876516, 6876553, 7939895, 6876554, 
    6876556, 11239240, 9640276, 789022, 789023, 6876559, 6876560, 7732816, 
    789024, 9977035, 10253225, 13596008, 13596009, 6876563, 6876562, 7732817, 
    6876564, 13596010, 6876567, 6876566, 7732818, 789027, 6876565, 789028, 
    6876523, 789025, 6876591, 9966446, 6876570, 789029, 7732819, 7506023, 
    6876577, 6876576, 6876574, 789030, 7939896, 789032, 6876573, 9977036, 
    9640277, 789034, 6876532, 789033, 6876579, 7732820, 7732821, 789036, 
    789035, 6876584, 6876580, 6876583, 9966447, 10253226, 9640278, 789037, 
    789039, 789040, 6876586, 789038, 6876546, 9977037, 789041, 789043, 
    7506024, 7939897, 789042, 11083086, 9640279, 789044, 6876589, 6876590, 
    6876598, 6876599, 6876596, 6876601, 6876600, 6876594, 789045, 6876593, 
    6876595, 6876597, 6876592 ;

 originators_station_identifier =
  "  ",
  "  ",
  "  ",
  "  ",
  "  ",
  "554_19,",
  "       ",
  "       ",
  "       ",
  "       ",
  "CWWSP",
  "     ",
  "     ",
  "     ",
  "     ",
  "     ",
  "     ",
  "     ",
  "     ",
  "     ",
  "     ",
  "     ",
  "     ",
  "     ",
  "     ",
  "     ",
  "     ",
  "     ",
  "     ",
  "     ",
  "     ",
  "     ",
  "     ",
  "     ",
  "     ",
  "     ",
  "     ",
  "     ",
  "     ",
  "     ",
  "     ",
  "     ",
  "     ",
  "554_20,",
  "       ",
  "TV",
  "TV",
  "  ",
  "  ",
  "  ",
  "  ",
  "TV",
  "  ",
  "  ",
  "  ",
  "  ",
  "  ",
  "  ",
  "  ",
  "  ",
  "  ",
  "  ",
  "  ",
  "  ",
  "  ",
  "  ",
  "  ",
  "  ",
  "  ",
  "  ",
  "  ",
  "  ",
  "  ",
  "  ",
  "  ",
  "  ",
  "  ",
  "  ",
  "  ",
  "  ",
  "  ",
  "  ",
  "  ",
  "  ",
  "  ",
  "  ",
  "  ",
  "  ",
  "  ",
  "  ",
  "  ",
  "  ",
  "  ",
  "  ",
  "  ",
  "  ",
  "554_21,",
  "       ",
  "       ",
  "       ",
  "       ",
  "       ",
  "       ",
  "       ",
  "       ",
  "       ",
  "       ",
  "       ",
  "       ",
  "       ",
  "       ",
  "       ",
  "       ",
  "       ",
  "       ",
  "       ",
  "       ",
  "       ",
  "       ",
  "       ",
  "       ",
  "       ",
  "       ",
  "       ",
  "       ",
  "       ",
  "       ",
  "       ",
  "       ",
  "       ",
  "       ",
  "       ",
  "       ",
  "       ",
  "       ",
  "       ",
  "       ",
  "       ",
  "       ",
  "554_22,",
  "       ",
  "       ",
  "       ",
  "       ",
  "       ",
  "       ",
  "       ",
  "       ",
  "       ",
  "       ",
  "       ",
  "       ",
  "       ",
  "       ",
  "       ",
  "       ",
  "       ",
  "       ",
  "       ",
  "       ",
  "TV",
  "  ",
  "  ",
  "  ",
  "  ",
  "  ",
  "  ",
  "  ",
  "  " ;

 lat = 26.68333, 3.15, 44.25, 40.51667, 40.817, 70.15, 57.93333, 34.96833, 
    43.55, 43.55, 71.50667, 42.03333, 44.13334, 57.85, 34.96833, 9, 36.46, 
    44.075, 40.233, 36, 34.96833, 71.25, 43.76667, 40.23333, 28.5, -0.33, 
    43.88334, 57.7, 20, 57.8, 40.71667, 34.87, 34.91833, 40.717, 57.63334, 
    34.81833, 34.86666, 56.28, 43.83333, 27.13333, 2.633333, 58.4, 43.6, 
    70.18333, 60.41667, 60.4, 58.38334, 43.76667, 8, -0.85, 36.63, 60.41667, 
    40.46667, 39.85, 57.7, 43.89167, 39.85, 70.99667, 20.03333, 58.33333, 
    40.467, 60.45, 60.43333, 29, 66.8, 58.26667, 43.43333, 43.95, -4.821667, 
    -24.27, 60.45, 51.175, 58.2, 60.46667, 44.08333, 34.51667, 43.33333, 
    40.31667, 40.21667, -18.43733, 57.9, 40.217, 40.317, 60.5, 27.61667, 
    58.13334, 11.31667, 56.6, 36.8, 43.36666, 16.05, -40.5, 57.81667, 
    51.12217, 44.15, 29.5, 70.16666, 39.75, 39.75, 70.74834, 58, 51.25, 20, 
    39.75, 57.63334, 70.505, 51.18616, 6.983334, -18.503, 44.26667, 40.567, 
    36, 40.56667, 35.06667, 57.93333, 44.4, 51.26117, 40.583, -18.552, 
    70.39833, 57.85, 43.73333, 28.06667, 40.58333, -40.5, 30, 37.3, 44.2, 
    40.733, 40.73333, 57.76667, 51.41667, 51.32784, 30.42333, 43.9, 20, 
    -18.58633, 57.7, 35.4, 70, 37.2, 44.325, 40.81667, 43.96667, -18.61867, 
    44.475, 40.817, 30.5, 44.58333, 44.70833, 41.067, 28.58333, 44.08333, 
    36.5, 37.03, 41.06667, 70.00333, 20, 53.33333, 53.16667, -28.76667, 
    53.33333, 40.22, 53.16667, 50, 53.33333, 53.33333, 53.33333, 53.33333 ;

 lon = 168.0167, 108.3667, -66.605, -71.6, -72.133, 56.33333, 9.45, 139.5533, 
    -59.86666, -59.8667, 31.22667, 153, -66.73333, 9.566667, 139.4667, -30, 
    -122.78, -66.61667, -71.95, -40, 139.3717, 31.215, -59.96667, -71.95, 
    141, -166.93, -66.63333, 9.783334, 137, 9.666667, -72.66666, 139.4367, 
    139.405, -72.667, 9.983334, 139.4683, -129.4333, -37, -66.46667, 169, 
    107.3833, 8.766666, -60.33333, 56.45, -1.35, -1.383333, 8.816667, 
    -66.41666, -30, -167.02, -122.38, -1.35, -73.21667, -72.45, 9.983334, 
    -66.28333, -72.45, 31.23167, 136, 8.9, -73.217, -1.316667, -1.333333, 
    141, 1.6, 8.983334, -60.58333, -66.425, 11.83833, 4.67, -1.3, 2.675, 
    9.083333, -1.316667, -66.43333, -130.1667, -60.75, -72.71667, -72.65, 
    36.97267, 10.45, -72.65, -72.717, -1.3, 169.9833, 9.183333, -32.71667, 
    -36.7, -122.07, -60.93333, -20.01667, -79.23333, 10.53333, 2.5055, 
    -66.38333, 141, 56.48333, 49.58333, 49.6, 31.21833, 9.366667, 2.616667, 
    134.9833, 49.61666, 10.71667, 31.21167, 2.452833, -30.01667, 37.13533, 
    -66.25, -72.467, -42.5, -72.46667, -130.6667, 9.466666, -66.13333, 
    2.3945, -72.45, 37.254, 31.21333, 9.566667, -60.63334, 170.95, -72.45, 
    -79.63333, 141, -122.62, -66.48333, -72.667, -72.66666, 9.7, 2.483333, 
    2.561167, -80.22, -61.05, 134, 37.33733, 9.75, -129.95, 56.06667, 
    -122.83, -66.34167, -72.13333, -61.41667, 37.41967, -66.24167, -72.133, 
    141, -66.11667, -65.98333, -71.7, 171.95, -61.25, 135.58, -123.2, -71.7, 
    30.61167, 133, 4, 4.483333, 114.3833, 3.266667, -72.65, 4.233333, -145, 
    4.5, 3.533333, 3.75, 4.25 ;

 time = 76769.0277778301, 76769, 76769.0291666668, 76769.0166666675, 
    76769.0374999978, 76769, 76769.0416666679, 76769.0791666657, 
    76769.0749999955, 76769.0756944418, 76769.0416666679, 76769.0625, 
    76769.0916666687, 76769.0854166672, 76769.1055555567, 76769.0833333358, 
    76769.140972212, 76769.1291666627, 76769.1379166692, 76769.125, 
    76769.1305555552, 76769.1458333284, 76769.1625000089, 76769.1416666657, 
    76769.125, 76769.125, 76769.200000003, 76769.2048611045, 
    76769.1666666716, 76769.1666666716, 76769.174999997, 76769.1958333254, 
    76769.1763888747, 76769.1716666669, 76769.2326388955, 76769.2194444537, 
    76769.211805582, 76769.2083333284, 76769.2666666806, 76769.2534722388, 
    76769.25, 76769.25, 76769.287499994, 76769.25, 76769.2916666567, 
    76769.2916666567, 76769.2916666567, 76769.3041666746, 76769.2916666567, 
    76769.2916666567, 76769.3715277612, 76769.3333333433, 76769.337500006, 
    76769.3583333492, 76769.34375, 76769.3666666746, 76769.349999994, 
    76769.3430555761, 76769.3333333433, 76769.3333333433, 76769.337500006, 
    76769.3333333433, 76769.3333333433, 76769.3333333433, 76769.375, 
    76769.375, 76769.3958333433, 76769.400000006, 76769.4458333254, 
    76769.4479166567, 76769.4166666567, 76769.4534722269, 76769.4166666567, 
    76769.4166666567, 76769.4541666508, 76769.4444444478, 76769.474999994, 
    76769.4874999821, 76769.4874999821, 76769.4715277851, 76769.46875, 
    76769.4779166877, 76769.4770833254, 76769.4583333433, 76769.4826388657, 
    76769.4583333433, 76769.4583333433, 76769.4583333433, 76769.5159721971, 
    76769.5374999642, 76769.5, 76769.5, 76769.5236111283, 76769.5, 
    76769.5333333611, 76769.5, 76769.5, 76769.511805594, 76769.5361111164, 
    76769.5534722209, 76769.5416666865, 76769.5500000119, 76769.5416666865, 
    76769.5534722209, 76769.6187500358, 76769.6201388836, 76769.59375, 
    76769.5833333135, 76769.5833333135, 76769.5875000358, 76769.5999999642, 
    76769.5833333135, 76769.6083333492, 76769.600694418, 76769.625, 
    76769.6374999881, 76769.625, 76769.6733333468, 76769.6666666865, 
    76769.6687499881, 76769.6666666865, 76769.679166615, 76769.6993055344, 
    76769.6708333492, 76769.6666666865, 76769.6666666865, 76769.7305555344, 
    76769.7458333373, 76769.7274999619, 76769.7375000119, 76769.7083333135, 
    76769.7173611522, 76769.7652778029, 76769.75, 76769.7791666985, 76769.75, 
    76769.75, 76769.75, 76769.7881944776, 76769.7534722686, 76769.8076388836, 
    76769.7916666865, 76769.8625000119, 76769.866666615, 76769.8333333135, 
    76769.8499999642, 76769.852083385, 76769.8333333135, 76769.9000000358, 
    76769.9541666508, 76769.9479166865, 76769.929166615, 76769.945833385, 
    76769.9166666865, 76769.9618055224, 76769.9875000119, 76769.9812499881, 
    76769.9583333135, 76769, 76769, 76769, 76769, 76769, 76769, 76769, 76769, 
    76769, 76769, 76769 ;

 date = 19800310, 19800310, 19800310, 19800310, 19800310, 19800310, 19800310, 
    19800310, 19800310, 19800310, 19800310, 19800310, 19800310, 19800310, 
    19800310, 19800310, 19800310, 19800310, 19800310, 19800310, 19800310, 
    19800310, 19800310, 19800310, 19800310, 19800310, 19800310, 19800310, 
    19800310, 19800310, 19800310, 19800310, 19800310, 19800310, 19800310, 
    19800310, 19800310, 19800310, 19800310, 19800310, 19800310, 19800310, 
    19800310, 19800310, 19800310, 19800310, 19800310, 19800310, 19800310, 
    19800310, 19800310, 19800310, 19800310, 19800310, 19800310, 19800310, 
    19800310, 19800310, 19800310, 19800310, 19800310, 19800310, 19800310, 
    19800310, 19800310, 19800310, 19800310, 19800310, 19800310, 19800310, 
    19800310, 19800310, 19800310, 19800310, 19800310, 19800310, 19800310, 
    19800310, 19800310, 19800310, 19800310, 19800310, 19800310, 19800310, 
    19800310, 19800310, 19800310, 19800310, 19800310, 19800310, 19800310, 
    19800310, 19800310, 19800310, 19800310, 19800310, 19800310, 19800310, 
    19800310, 19800310, 19800310, 19800310, 19800310, 19800310, 19800310, 
    19800310, 19800310, 19800310, 19800310, 19800310, 19800310, 19800310, 
    19800310, 19800310, 19800310, 19800310, 19800310, 19800310, 19800310, 
    19800310, 19800310, 19800310, 19800310, 19800310, 19800310, 19800310, 
    19800310, 19800310, 19800310, 19800310, 19800310, 19800310, 19800310, 
    19800310, 19800310, 19800310, 19800310, 19800310, 19800310, 19800310, 
    19800310, 19800310, 19800310, 19800310, 19800310, 19800310, 19800310, 
    19800310, 19800310, 19800310, 19800310, 19800310, 19800310, 19800310, 
    19800310, 19800310, 19800310, 19800310, 19800310, 19800310, 19800310, 
    19800310, 19800310, 19800310, 19800310, 19800310, 19800310, 19800310, 
    19800310 ;

 GMT_time = 0.6666679, 0, 0.7, 0.4, 0.9, 0, 1, 1.9, 1.8, 1.816667, 1, 1.5, 
    2.2, 2.05, 2.533333, 2, 3.383333, 3.1, 3.31, 3, 3.133333, 3.5, 3.9, 3.4, 
    3, 3, 4.8, 4.916667, 4, 4, 4.2, 4.7, 4.233333, 4.12, 5.583333, 5.266667, 
    5.083334, 5, 6.4, 6.083334, 6, 6, 6.9, 6, 7, 7, 7, 7.3, 7, 7, 8.916666, 
    8, 8.1, 8.6, 8.25, 8.8, 8.4, 8.233334, 8, 8, 8.1, 8, 8, 8, 9, 9, 9.5, 
    9.6, 10.7, 10.75, 10, 10.88333, 10, 10, 10.9, 10.66667, 11.4, 11.7, 11.7, 
    11.31667, 11.25, 11.47, 11.45, 11, 11.58333, 11, 11, 11, 12.38333, 12.9, 
    12, 12, 12.56667, 12, 12.8, 12, 12, 12.28333, 12.86667, 13.28333, 13, 
    13.2, 13, 13.28333, 14.85, 14.88333, 14.25, 14, 14, 14.1, 14.4, 14, 14.6, 
    14.41667, 15, 15.3, 15, 16.16, 16, 16.05, 16, 16.3, 16.78333, 16.1, 16, 
    16, 17.53333, 17.9, 17.46, 17.7, 17, 17.21667, 18.36667, 18, 18.7, 18, 
    18, 18, 18.91667, 18.08333, 19.38333, 19, 20.7, 20.8, 20, 20.4, 20.45, 
    20, 21.6, 22.9, 22.75, 22.3, 22.7, 22, 23.08333, 23.7, 23.55, 23, _, _, 
    _, _, _, _, _, _, _, _, _ ;

 Access_no = 273, 8300094, 8200231, 8100661, 2023, 71066, 9600121, 416, 
    8200231, 9600170, 9600121, 526, 8200231, 9600121, 416, 8300094, 1021, 
    8200231, 9800126, 8300094, 416, 9600121, 8200231, 8100661, 937, 38350, 
    8200231, 9600121, 9700253, 9600121, 204, 416, 416, 9800126, 9600121, 416, 
    526, 38350, 8200231, 273, 8300094, 9500146, 8200231, 71066, 9700138, 
    9700138, 9500146, 8200231, 8300094, 38350, 1021, 9700138, 204, 8100661, 
    9600121, 8200231, 9800126, 9600121, 9700253, 9600121, 9800126, 9700138, 
    9700138, 937, 9700164, 9600121, 8200231, 8200231, 8600187, 305, 9700138, 
    101, 9600121, 9700138, 8200231, 526, 8200231, 204, 8100661, 9200135, 
    9600121, 9800126, 9800126, 9700138, 273, 9600121, 9700253, 38350, 1021, 
    8200231, 8300094, 9700249, 9600121, 101, 8200231, 937, 71066, 72200, 
    72200, 9600121, 9600121, 101, 9700253, 72200, 9600121, 9600121, 101, 
    8300094, 9200135, 8200231, 9800126, 8300094, 204, 526, 9600121, 8200231, 
    101, 9800126, 9200135, 9600121, 9600121, 8200231, 273, 8100661, 9700249, 
    937, 1021, 8200231, 9800126, 8100661, 9600121, 101, 101, 8500245, 
    8200231, 9700253, 9200135, 9600121, 526, 71066, 1021, 8200231, 8100661, 
    8200231, 9200135, 8200231, 9800126, 937, 8200231, 8200231, 9800126, 273, 
    8200231, 31246, 1021, 8100661, 9600121, 9700253, 9700138, 9700138, 
    9200118, 9700138, 9400135, 9700138, 8900177, 9700138, 9700138, 9700138, 
    9700138 ;

 Project =
  "MARINE RESOURCES MONITORING ASSESSMENT & PREDICTION PROGRAM (MARMAP)",
  "POD (1963 - 1996)",
  "POD (1963 - 1996)",
  "MARINE RESOURCES MONITORING ASSESSMENT & PREDICTION PROGRAM (MARMAP)",
  "POD (1963 - 1996)",
  "MARINE RESOURCES MONITORING ASSESSMENT & PREDICTION PROGRAM (MARMAP)",
  "MARINE RESOURCES MONITORING ASSESSMENT & PREDICTION PROGRAM (MARMAP)",
  "POD (1963 - 1996)",
  "POD (1963 - 1996)",
  "MARINE RESOURCES MONITORING ASSESSMENT & PREDICTION PROGRAM (MARMAP)",
  "POD (1963 - 1996)",
  "MARINE RESOURCES MONITORING ASSESSMENT & PREDICTION PROGRAM (MARMAP)",
  "MARINE RESOURCES MONITORING ASSESSMENT & PREDICTION PROGRAM (MARMAP)",
  "MARINE RESOURCES MONITORING ASSESSMENT & PREDICTION PROGRAM (MARMAP)",
  "MARINE RESOURCES MONITORING ASSESSMENT & PREDICTION PROGRAM (MARMAP)",
  "MARINE RESOURCES MONITORING ASSESSMENT & PREDICTION PROGRAM (MARMAP)",
  "MARINE RESOURCES MONITORING ASSESSMENT & PREDICTION PROGRAM (MARMAP)",
  "MARINE RESOURCES MONITORING ASSESSMENT & PREDICTION PROGRAM (MARMAP)",
  "MARINE RESOURCES MONITORING ASSESSMENT & PREDICTION PROGRAM (MARMAP)",
  "MARINE RESOURCES MONITORING ASSESSMENT & PREDICTION PROGRAM (MARMAP)",
  "MARINE RESOURCES MONITORING ASSESSMENT & PREDICTION PROGRAM (MARMAP)",
  "MARINE RESOURCES MONITORING ASSESSMENT & PREDICTION PROGRAM (MARMAP)",
  "MARINE RESOURCES MONITORING ASSESSMENT & PREDICTION PROGRAM (MARMAP)",
  "MARINE RESOURCES MONITORING ASSESSMENT & PREDICTION PROGRAM (MARMAP)",
  "MARINE RESOURCES MONITORING ASSESSMENT & PREDICTION PROGRAM (MARMAP)",
  "MARINE RESOURCES MONITORING ASSESSMENT & PREDICTION PROGRAM (MARMAP)",
  "MARINE RESOURCES MONITORING ASSESSMENT & PREDICTION PROGRAM (MARMAP)",
  "MARINE RESOURCES MONITORING ASSESSMENT & PREDICTION PROGRAM (MARMAP)",
  "MARINE RESOURCES MONITORING ASSESSMENT & PREDICTION PROGRAM (MARMAP)",
  "MARINE RESOURCES MONITORING ASSESSMENT & PREDICTION PROGRAM (MARMAP)",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "" ;

 Platform =
  "SHOYO MARU",
  "AKADEMIK KOROLYOV (R/V; call sign UHQS; built 06.1967; IMO6707301)",
  "E. E. PRINCE (AFTER 1960)",
  "ALBATROSS IV (NOAA ship; call sign WMVF; built 1962; IMO7338690)",
  "WIECZNO",
  "OTTO SCHMIDT (1979)",
  "JOHAN HJORT (R/V;call sign LDGJ; built 1990; IMO8915768)!",
  "USHIO (Built 01.1991)",
  "LADY HAMMOND",
  "A. T. CAMERON",
  "G.O. SARS (R/V; call sign LLZG; active 1970-2003;IMO7018379)",
  "MYS DALNIY (F/V; call sign UWKC; built 1977; IMO7643942)!",
  "E. E. PRINCE (AFTER 1960)",
  "JOHAN HJORT (R/V;call sign LDGJ; built 1990; IMO8915768)!",
  "USHIO (Built 01.1991)",
  "ERNST KRENKEL (R/V;c.s.EREU;built1971;ex.Vikhr 1972;n.c.s.EOGQ;IMO7205685)",
  "TIKHOOKEANSKIY (Call sign EUEM; built 1976; IMO7640897)",
  "E. E. PRINCE (AFTER 1960)",
  "ALBATROSS IV (NOAA ship; call sign WMVF; built 1962; IMO7338690)",
  "MUSSON (R/V; call sign EREA; built 1968; decomm-d 1992;IMO6904155)",
  "USHIO (Built 01.1991)",
  "G.O. SARS (R/V; call sign LLZG; active 1970-2003;IMO7018379)",
  "LADY HAMMOND",
  "ALBATROSS IV (NOAA ship; call sign WMVF; built 1962; IMO7338690)",
  "VOLNA",
  "DMITRIY MENDELEYEV (R/V; call sign UILS; built 1968; IMO6806896)",
  "E. E. PRINCE (AFTER 1960)",
  "JOHAN HJORT (R/V;call sign LDGJ; built 1990; IMO8915768)!",
  "OKEAN",
  "JOHAN HJORT (R/V;call sign LDGJ; built 1990; IMO8915768)!",
  "WIECZNO",
  "USHIO (Built 01.1991)",
  "USHIO (Built 01.1991)",
  "WIECZNO",
  "JOHAN HJORT (R/V;call sign LDGJ; built 1990; IMO8915768)!",
  "USHIO (Built 01.1991)",
  "NOVOULYANOVSK (R/V; call sign UKGF; built 1979; IMO7932757)",
  "AYAKS (F/V; call sign UUWI; built 1972; IMO7304194; Murmansk)",
  "E. E. PRINCE (AFTER 1960)",
  "SHOYO MARU",
  "AKADEMIK KOROLYOV (R/V; call sign UHQS; built 06.1967; IMO6707301)",
  "LADY HAMMOND",
  "OTTO SCHMIDT (1979)",
  "MARA",
  "MARA",
  "E. E. PRINCE (AFTER 1960)",
  "ERNST KRENKEL (R/V;c.s.EREU;built1971;ex.Vikhr 1972;n.c.s.EOGQ;IMO7205685)",
  "DMITRIY MENDELEYEV (R/V; call sign UILS; built 1968; IMO6806896)",
  "TIKHOOKEANSKIY (Call sign EUEM; built 1976; IMO7640897)",
  "MARA",
  "WIECZNO",
  "ALBATROSS IV (NOAA ship; call sign WMVF; built 1962; IMO7338690)",
  "JOHAN HJORT (R/V;call sign LDGJ; built 1990; IMO8915768)!",
  "E. E. PRINCE (AFTER 1960)",
  "ALBATROSS IV (NOAA ship; call sign WMVF; built 1962; IMO7338690)",
  "G.O. SARS (R/V; call sign LLZG; active 1970-2003;IMO7018379)",
  "OKEAN",
  "G.M. DANNEVIG (R/V;call sign LINW;built 1979;ex.Kystfangst 1987;IMO8899665)",
  "WIECZNO",
  "MARA",
  "MARA",
  "VOLNA",
  "G.M. DANNEVIG (R/V;call sign LINW;built 1979;ex.Kystfangst 1987;IMO8899665)",
  "LADY HAMMOND",
  "E. E. PRINCE (AFTER 1960)",
  "WHARF POINTE NOIRE",
  "60 LET VLKSM (F/V; call sign EWYB; built 1978; IMO 7740776; Zapryba)",
  "MARA",
  "MECHELEN",
  "G.M. DANNEVIG (R/V;call sign LINW;built 1979;ex.Kystfangst 1987;IMO8899665)",
  "MARA",
  "E. E. PRINCE (AFTER 1960)",
  "NOVOULYANOVSK (R/V; call sign UKGF; built 1979; IMO7932757)",
  "LADY HAMMOND",
  "WIECZNO",
  "ALBATROSS IV (NOAA ship; call sign WMVF; built 1962; IMO7338690)",
  "A.V.HUMBOLDT (R/V;c.s.Y3CW;comm-d 1970;decomm-d 1990;IMO6711883)",
  "JOHAN HJORT (R/V;call sign LDGJ; built 1990; IMO8915768)!",
  "ALBATROSS IV (NOAA ship; call sign WMVF; built 1962; IMO7338690)",
  "WIECZNO",
  "MARA",
  "SHOYO MARU",
  "G.M. DANNEVIG (R/V;call sign LINW;built 1979;ex.Kystfangst 1987;IMO8899665)",
  "SRTM 8005 \"ALIOT\"",
  "AYAKS (F/V; call sign UUWI; built 1972; IMO7304194; Murmansk)",
  "TIKHOOKEANSKIY (Call sign EUEM; built 1976; IMO7640897)",
  "LADY HAMMOND",
  "PASSAT (R/V;c.s.UZGH;b.1968;IMOO6904167;flag USSR; Ukraine 1993-2008)",
  "ZVEZDA KRIMA (R/F/V; call sign UWGM; built 1972; IMO7229526)",
  "JOHAN HJORT (R/V;call sign LDGJ; built 1990; IMO8915768)!",
  "MECHELEN",
  "E. E. PRINCE (AFTER 1960)",
  "VOLNA",
  "OTTO SCHMIDT (1979)",
  "OKEANOLOG (Small boat)",
  "OKEANOLOG (Small boat)",
  "G.O. SARS (R/V; call sign LLZG; active 1970-2003;IMO7018379)",
  "G.M. DANNEVIG (R/V;call sign LINW;built 1979;ex.Kystfangst 1987;IMO8899665)",
  "MECHELEN",
  "OKEAN",
  "OKEANOLOG (Small boat)",
  "JOHAN HJORT (R/V;call sign LDGJ; built 1990; IMO8915768)!",
  "G.O. SARS (R/V; call sign LLZG; active 1970-2003;IMO7018379)",
  "MECHELEN",
  "ERNST KRENKEL (R/V;c.s.EREU;built1971;ex.Vikhr 1972;n.c.s.EOGQ;IMO7205685)",
  "A.V.HUMBOLDT (R/V;c.s.Y3CW;comm-d 1970;decomm-d 1990;IMO6711883)",
  "E. E. PRINCE (AFTER 1960)",
  "WIECZNO",
  "MUSSON (R/V; call sign EREA; built 1968; decomm-d 1992;IMO6904155)",
  "WIECZNO",
  "NOVOULYANOVSK (R/V; call sign UKGF; built 1979; IMO7932757)",
  "G.M. DANNEVIG (R/V;call sign LINW;built 1979;ex.Kystfangst 1987;IMO8899665)",
  "E. E. PRINCE (AFTER 1960)",
  "MECHELEN",
  "ALBATROSS IV (NOAA ship; call sign WMVF; built 1962; IMO7338690)",
  "A.V.HUMBOLDT (R/V;c.s.Y3CW;comm-d 1970;decomm-d 1990;IMO6711883)",
  "G.O. SARS (R/V; call sign LLZG; active 1970-2003;IMO7018379)",
  "G.M. DANNEVIG (R/V;call sign LINW;built 1979;ex.Kystfangst 1987;IMO8899665)",
  "LADY HAMMOND",
  "SHOYO MARU",
  "ALBATROSS IV (NOAA ship; call sign WMVF; built 1962; IMO7338690)",
  "ZVEZDA KRIMA (R/F/V; call sign UWGM; built 1972; IMO7229526)",
  "VOLNA",
  "TIKHOOKEANSKIY (Call sign EUEM; built 1976; IMO7640897)",
  "E. E. PRINCE (AFTER 1960)",
  "ALBATROSS IV (NOAA ship; call sign WMVF; built 1962; IMO7338690)",
  "ALBATROSS IV (NOAA ship; call sign WMVF; built 1962; IMO7338690)",
  "G.M. DANNEVIG (R/V;call sign LINW;built 1979;ex.Kystfangst 1987;IMO8899665)",
  "MECHELEN",
  "MECHELEN",
  "DARBY",
  "LADY HAMMOND",
  "OKEAN",
  "A.V.HUMBOLDT (R/V;c.s.Y3CW;comm-d 1970;decomm-d 1990;IMO6711883)",
  "G.M. DANNEVIG (R/V;call sign LINW;built 1979;ex.Kystfangst 1987;IMO8899665)",
  "NOVOULYANOVSK (R/V; call sign UKGF; built 1979; IMO7932757)",
  "OTTO SCHMIDT (1979)",
  "TIKHOOKEANSKIY (Call sign EUEM; built 1976; IMO7640897)",
  "E. E. PRINCE (AFTER 1960)",
  "ALBATROSS IV (NOAA ship; call sign WMVF; built 1962; IMO7338690)",
  "LADY HAMMOND",
  "A.V.HUMBOLDT (R/V;c.s.Y3CW;comm-d 1970;decomm-d 1990;IMO6711883)",
  "E. E. PRINCE (AFTER 1960)",
  "ALBATROSS IV (NOAA ship; call sign WMVF; built 1962; IMO7338690)",
  "VOLNA",
  "E. E. PRINCE (AFTER 1960)",
  "E. E. PRINCE (AFTER 1960)",
  "ALBATROSS IV (NOAA ship; call sign WMVF; built 1962; IMO7338690)",
  "SHOYO MARU",
  "LADY HAMMOND",
  "PRIBOY",
  "TIKHOOKEANSKIY (Call sign EUEM; built 1976; IMO7640897)",
  "ALBATROSS IV (NOAA ship; call sign WMVF; built 1962; IMO7338690)",
  "G.O. SARS (R/V; call sign LLZG; active 1970-2003;IMO7018379)",
  "OKEAN",
  "CIROLANA",
  "CIROLANA",
  "GERALDTON",
  "CIROLANA",
  "CIROLANA",
  "VANCOUVER (Old OWS \'P\' reporting vessel)!",
  "CIROLANA",
  "CIROLANA",
  "CIROLANA",
  "CIROLANA",
  "",
  "",
  "",
  "" ;

 Institute =
  "FISHERIES AGENCY OF JAPAN (JFA) TOKYO",
  "HYDROMETEOROLOGICAL SERVICE (MOSCOW)",
  "US DOC NOAA NMFS (WOODS HOLE; MA)",
  "ARCTIC AND ANTARCTIC RESEARCH INSTITUTE (AARI)",
  "SAGAMI BAY EXPERIMENTAL STATION",
  "PACIFIC RES INST OF FISH AND OCY (TINRO; AND OTHERS)",
  "SAGAMI BAY EXPERIMENTAL STATION",
  "HYDROMETEOROLOGICAL SERVICE (MOSCOW)",
  "PACIFIC RES INST OF FISH AND OCY (TINRO; AND OTHERS)",
  "US DOC NOAA NMFS (NARRAGANSETT; RI)",
  "HYDROMETEOROLOGICAL SERVICE (MOSCOW)",
  "SAGAMI BAY EXPERIMENTAL STATION",
  "US DOC NOAA NMFS (WOODS HOLE; MA)",
  "FAR EASTERN REGIONAL HYDROMETEOROLOGICAL RESEARCH INSTITUTE; FERHRI",
  "P.P.SHIRSHOV INSTITUTE OF OCEANOLOGY OF THE RUSSIAN ACADEMY OF SCIENCES",
  "FAR EASTERN REGIONAL HYDROMETEOROLOGICAL RESEARCH INSTITUTE; FERHRI",
  "SAGAMI BAY EXPERIMENTAL STATION",
  "SAGAMI BAY EXPERIMENTAL STATION",
  "US DOC NOAA NMFS (NARRAGANSETT; RI)",
  "SAGAMI BAY EXPERIMENTAL STATION",
  "PACIFIC RES INST OF FISH AND OCY (TINRO; AND OTHERS)",
  "POLAR RES AND DESIGNING INST OF MARINE FISH AND OCY PINRO (MURMANSK)",
  "FISHERIES AGENCY OF JAPAN (JFA) TOKYO",
  "HYDROMETEOROLOGICAL SERVICE (MOSCOW)",
  "ARCTIC AND ANTARCTIC RESEARCH INSTITUTE (AARI)",
  "HYDROMETEOROLOGICAL SERVICE (MOSCOW)",
  "P.P.SHIRSHOV INSTITUTE OF OCEANOLOGY OF THE RUSSIAN ACADEMY OF SCIENCES",
  "PACIFIC RES INST OF FISH AND OCY (TINRO; AND OTHERS)",
  "US DOC NOAA NMFS (WOODS HOLE; MA)",
  "US DOC NOAA NMFS (NARRAGANSETT; RI)",
  "FAR EASTERN REGIONAL HYDROMETEOROLOGICAL RESEARCH INSTITUTE; FERHRI",
  "US DOC NOAA NMFS (NARRAGANSETT; RI)",
  "FAR EASTERN REGIONAL HYDROMETEOROLOGICAL RESEARCH INSTITUTE; FERHRI",
  "CENTRE NATIONAL POUR L\'EXPLOITATION DES OCEANS (CNEXO)",
  "ATLANTIC RESEARCH INST OF FISHING ECONOMY AND OCEANOGRAPHY (ATLANTNIRO)",
  "PACIFIC RES INST OF FISH AND OCY (TINRO; AND OTHERS)",
  "US DOC NOAA NMFS (WOODS HOLE; MA)",
  "US DOC NOAA NMFS (NARRAGANSETT; RI)",
  "US DOC NOAA NMFS (NARRAGANSETT; RI)",
  "FISHERIES AGENCY OF JAPAN (JFA) TOKYO",
  "ATLANTIC RESEARCH INST OF FISHING ECONOMY AND OCEANOGRAPHY (ATLANTNIRO)",
  "POLAR RES AND DESIGNING INST OF MARINE FISH AND OCY PINRO (MURMANSK)",
  "PACIFIC RES INST OF FISH AND OCY (TINRO; AND OTHERS)",
  "HYDROMETEOROLOGICAL SERVICE (MOSCOW)",
  "FAR EASTERN REGIONAL HYDROMETEOROLOGICAL RESEARCH INSTITUTE; FERHRI",
  "ARCTIC AND ANTARCTIC RESEARCH INSTITUTE (AARI)",
  "HYDROMETEOROLOGICAL SERVICE (AZERBAJAN)",
  "HYDROMETEOROLOGICAL SERVICE (AZERBAJAN)",
  "FAR EASTERN REGIONAL HYDROMETEOROLOGICAL RESEARCH INSTITUTE; FERHRI",
  "HYDROMETEOROLOGICAL SERVICE (AZERBAJAN)",
  "HYDROMETEOROLOGICAL SERVICE (MOSCOW)",
  "US DOC NOAA NMFS (NARRAGANSETT; RI)",
  "HYDROMETEOROLOGICAL SERVICE (MOSCOW)",
  "PACIFIC RES INST OF FISH AND OCY (TINRO; AND OTHERS)",
  "US DOC NOAA NMFS (NARRAGANSETT; RI)",
  "FISHERIES AGENCY OF JAPAN (JFA) TOKYO",
  "US DOC NOAA NMFS (WOODS HOLE; MA)",
  "FAR EASTERN REGIONAL HYDROMETEOROLOGICAL RESEARCH INSTITUTE; FERHRI",
  "PACIFIC RES INST OF FISH AND OCY (TINRO; AND OTHERS)",
  "US DOC NOAA NMFS (NARRAGANSETT; RI)",
  "US DOC NOAA NMFS (WOODS HOLE; MA)",
  "MARINE RESOURCES RESEARCH INST (CHARLESTON; SC)",
  "FAR EASTERN REGIONAL HYDROMETEOROLOGICAL RESEARCH INSTITUTE; FERHRI",
  "PACIFIC RES INST OF FISH AND OCY (TINRO; AND OTHERS)",
  "ARCTIC AND ANTARCTIC RESEARCH INSTITUTE (AARI)",
  "PACIFIC RES INST OF FISH AND OCY (TINRO; AND OTHERS)",
  "US DOC NOAA NMFS (WOODS HOLE; MA)",
  "US DOC NOAA NMFS (NARRAGANSETT; RI)",
  "FAR EASTERN REGIONAL HYDROMETEOROLOGICAL RESEARCH INSTITUTE; FERHRI",
  "US DOC NOAA NMFS (NARRAGANSETT; RI)",
  "FISHERIES AGENCY OF JAPAN (JFA) TOKYO",
  "FAR EASTERN REGIONAL HYDROMETEOROLOGICAL RESEARCH INSTITUTE; FERHRI",
  "PACIFIC RES INST OF FISH AND OCY (TINRO; AND OTHERS)",
  "US DOC NOAA NMFS (WOODS HOLE; MA)",
  "FAR EASTERN REGIONAL HYDROMETEOROLOGICAL RESEARCH INSTITUTE; FERHRI",
  "CANADIAN OCEANOGRAPHIC DATA CENTER (OTTAWA) ** USE CODE 1199 **",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "" ;

 Orig_Stat_Num = _, _, _, 67, _, _, _, _, _, 29, _, 109, _, _, _, _, 63, _, 
    68, _, _, _, _, 68, 123, 27, _, _, 39, _, 89, _, _, 89, _, _, 30, 26, _, 
    _, _, _, _, _, _, _, _, _, _, 28, 64, _, 90, 69, _, _, 69, _, 40, _, 90, 
    _, _, 124, _, _, _, _, _, 25, _, _, _, _, _, 31, _, 91, 70, _, _, 70, 91, 
    _, _, _, 34, 27, 65, _, _, 9500, _, _, _, 125, _, 1, 2, _, _, _, 41, 3, 
    _, _, _, _, _, _, 92, _, 92, 32, _, _, _, 71, _, _, _, _, _, 71, 9600, 
    126, 66, _, 72, 72, _, _, _, 3320365, _, 42, _, _, 33, _, 67, _, 73, _, 
    _, _, 73, 127, _, _, 74, _, _, 220, 68, 74, _, 43, _, _, _, _, _, _, 42, 
    _, _, _, _ ;

 Bottom_Depth = _, 80, 197, 73, 37, 110, _, _, 270, 270, _, 5280, 73, _, _, 
    5300, 3040, 95, _, 4000, _, _, 56, 66, 3800, 5800, 95, _, 4600, _, 32, _, 
    _, _, _, _, 4900, 2440, 65, _, 80, 110, 70, 105, 26, 36, 90, 84, 4470, 
    5820, 2750, 17, 28, 71, _, 36, _, _, 4700, 240, _, 23, 25, 3950, 2000, 
    400, 108, 69, 18, 3250, 17, _, 420, 17, 76, 4900, 277, 53, 57, 26, _, _, 
    _, 51, _, 640, 5800, 2600, 215, 109, 3600, 4100, _, _, 69, 3900, 105, 13, 
    12, _, 400, _, 5700, 11, _, _, _, 4170, 35, 38, _, 4260, 38, 4700, 190, 
    29, _, _, 83, _, 90, 53, _, 44, 4500, 3400, 87, 100, _, 26, 32, _, _, 59, 
    52, 4580, 350, 65, 4500, 85, 325, 76, 37, 75, 780, 95, _, 3100, 88, 95, 
    _, _, 87, _, 2300, 53, _, 6000, 30, 31, 40, 27, _, 31, _, 29, 28, 28, 28 ;

 Cast_Duration = _, _, _, _, _, _, _, _, _, _, _, 1.166667, _, _, _, _, _, _, 
    _, _, _, _, _, _, 1, _, _, _, _, _, _, _, _, _, _, _, 0.5833321, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 2, 
    _, _, _, _, _, 0.916667, _, _, _, _, _, 0.666666, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, 1, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, 0.5, _, _, _, _, _, _, _, _, _, _, _, 1, _, _, _, _, _, _, 
    _, _, _, _, _, _, 0.5833321, _, _, _, _, _, _, _, _, 2, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 Water_Color =
  "PERCENT YELLOW 5  FOREL-ULE SCALE III",
  "PERCENT YELLOW 5  FOREL-ULE SCALE III",
  "PERCENT YELLOW 5  FOREL-ULE SCALE III",
  "PERCENT YELLOW 5  FOREL-ULE SCALE III",
  "PERCENT YELLOW 5  FOREL-ULE SCALE III",
  "PERCENT YELLOW 35  FOREL-ULE SCALE VIII",
  "PERCENT YELLOW 35  FOREL-ULE SCALE VIII",
  "PERCENT YELLOW 35  FOREL-ULE SCALE VIII",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "" ;

 Water_Transpar = _, _, _, _, _, _, _, 2, _, _, _, _, _, _, _, _, _, _, _, _, 
    2, _, _, _, _, _, _, _, _, _, _, 2, 2, _, _, 2, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, 5, 5, _, _, _, _, 5, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _ ;

 Wave_Direction =
  "15 DEGREES - 24 DEGREES",
  "285 DEGREES - 294 DEGREES",
  "5 DEGREES - 14 DEGREES",
  "5 DEGREES - 14 DEGREES",
  "5 DEGREES - 14 DEGREES",
  "315 DEGREES - 324 DEGREES",
  "135 DEGREES - 144 DEGREES",
  "45 DEGREES - 54 DEGREES",
  "45 DEGREES - 54 DEGREES",
  "45 DEGREES - 54 DEGREES",
  "295 DEGREES - 304 DEGREES",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "" ;

 Wave_Height =
  "4 METER",
  "3 METER",
  "2.5 METER",
  "1.5 METER",
  "3.5 METER",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "" ;

 Sea_State =
  "CALM-GLASSY 0 FT (0 METERS)",
  "SLIGHT 1 2/3 - 4 FT(.5-1.25 METERS)",
  "VERY ROUGH 13-20 FT(4-6 METERS)",
  "SLIGHT 1 2/3 - 4 FT(.5-1.25 METERS)",
  "SLIGHT 1 2/3 - 4 FT(.5-1.25 METERS)",
  "CALM-RIPPLED 0-1/3 FT (0-.1METERS)",
  "VERY ROUGH 13-20 FT(4-6 METERS)",
  "MODERATE 4-8 FT(1.25-2.50 METERS)",
  "CALM-RIPPLED 0-1/3 FT (0-.1METERS)",
  "CALM MEAN VELOCITY IN KNOTS <1 IN METERS/SEC 0-0.2 IN KM/H <1 IN M.P.H. <1 /WAVE HT < .25 FT",
  "CALM MEAN VELOCITY IN KNOTS <1 IN METERS/SEC 0-0.2 IN KM/H <1 IN M.P.H. <1 /WAVE HT < .25 FT",
  "CALM MEAN VELOCITY IN KNOTS <1 IN METERS/SEC 0-0.2 IN KM/H <1 IN M.P.H. <1 /WAVE HT < .25 FT",
  "VERY ROUGH 13-20 FT(4-6 METERS)",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "" ;

 Wind_Force =
  "LIGHT AIR  MEAN VELOCITY IN KNOTS 1-3  METERS/SEC 0.3-1.5 KM/H 1-5 M.P.H. 1-3 /WAVE HT= .25 FT",
  "MODERATE BREEZE  MEAN VELOCITY IN KNOTS 11-16  METERS/SEC 5.5-7.9  KM/H 20-28  M.P.H. 13-18 WAVE HT = 4 FT",
  "GENTLE BREEZE  MEAN VELOCITY IN KNOTS 7-10  METERS/SEC 3.4-5.4  KM/H 12-19  M.P.H. 8-12 /WAVE HT = 2 FT",
  "MODERATE BREEZE  MEAN VELOCITY IN KNOTS 11-16  METERS/SEC 5.5-7.9  KM/H 20-28  M.P.H. 13-18 WAVE HT = 4 FT",
  "LIGHT BREEZE  MEAN VELOCITY IN KNOTS 4-6  METERS/SEC 1.6-3.3 KM/H 6-11  M.P.H. 4-7 /WAVE HT = .5 FT",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "" ;

 Wave_Period =
  "5 SECONDS OR LESS",
  "5 SECONDS OR LESS",
  "5 SECONDS OR LESS",
  "5 SECONDS OR LESS",
  "5 SECONDS OR LESS",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "" ;

 Wind_Direction =
  "235 DEGREES - 244 DEGREES",
  "85 DEGREES - 94 DEGREES",
  "145 DEGREES - 154 DEGREES",
  "285 DEGREES - 294 DEGREES",
  "105 DEGREES - 114 DEGREES",
  "85 DEGREES - 94 DEGREES",
  "105 DEGREES - 114 DEGREES",
  "45 DEGREES - 54 DEGREES",
  "225 DEGREES - 234 DEGREES",
  "315 DEGREES - 324 DEGREES",
  "135 DEGREES - 144 DEGREES",
  "45 DEGREES - 54 DEGREES",
  "315 DEGREES - 324 DEGREES",
  "225 DEGREES - 234 DEGREES",
  "45 DEGREES - 54 DEGREES",
  "45 DEGREES - 54 DEGREES",
  "45 DEGREES - 54 DEGREES",
  "45 DEGREES - 54 DEGREES",
  "295 DEGREES - 304 DEGREES",
  "355 DEGREES - 4 DEGREES",
  "CALM (NO WAVES-NO MOTION)",
  "215 DEGREES - 224 DEGREES",
  "295 DEGREES - 304 DEGREES",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "" ;

 Wind_Speed = _, _, _, _, _, 13.608, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, 31.104, _, _, _, _, _, _, _, _, _, _, _, 25.272, _, _, _, 
    _, _, _, 9.72, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    25.272, _, _, _, _, _, 19.8288, _, _, _, _, _, 21.384, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, 23.328, 11.664, 7.776, 7.776, _, 
    _, _, _, 7.776, _, _, _, _, _, _, _, _, _, 21.384, _, _, _, _, _, _, _, 
    _, _, _, _, 17.496, _, _, _, _, _, _, _, _, _, _, _, _, 16.3296, 13.608, 
    _, _, _, _, _, _, _, 23.328, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _ ;

 Barometric_Pres = _, _, _, _, _, 1035, _, 1000, _, _, _, _, _, _, _, _, _, 
    _, _, _, 1001, _, _, _, 1008.7, _, _, _, _, _, _, 1001.5, 1001, _, _, 
    1002.5, 1021.9, _, _, _, _, _, _, 1034.6, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, 1010.1, _, _, _, _, _, 1026.3, _, _, _, _, _, 
    1020.9, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 1011.3, 
    1034, 1026.9, 1026.8, _, _, _, _, 1026.8, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, 1011, _, _, _, _, _, _, _, 1013.2, _, _, 
    _, _, 1023, 1033.4, _, _, _, _, _, _, _, 1012.1, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 Dry_Bulb_Temp = _, _, _, _, _, -6.6, _, 15, _, _, _, _, _, _, _, _, _, _, _, 
    _, 17.5, _, _, _, 19.2, _, _, _, _, _, _, 17, 16.8, _, _, 17, 13.6, _, _, 
    _, _, _, _, -8.7, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, 17.6, _, _, _, _, _, 22.3, _, _, _, _, _, 13.6, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, 17.7, -6.6, 7.2, 7.1, _, _, _, _, 7, 
    _, _, _, _, _, _, _, _, _, 12.6, _, _, _, _, _, _, _, _, _, _, _, 15.7, 
    _, _, _, _, _, _, _, 19.4, _, _, _, _, 12.7, -11.6, _, _, _, _, _, _, _, 
    14.8, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 Weather_Condition =
  "STATE OF SKY ON THE WHOLE UNCHANGED-CHAR. CHANGE OF THE STATE OF SKY DURING THE PAST HOUR",
  "CLEAR (NO CLOUD AT ANY LEVEL)",
  "CLEAR (NO CLOUD AT ANY LEVEL)",
  "STATE OF SKY ON THE WHOLE UNCHANGED-CHAR. CHANGE OF THE STATE OF SKY DURING THE PAST HOUR",
  "CLEAR (NO CLOUD AT ANY LEVEL)",
  "CLEAR (NO CLOUD AT ANY LEVEL)",
  "CLEAR (NO CLOUD AT ANY LEVEL)",
  "CLOUDS GENERALLY DISSOLVING OF BECOMING LESS DEVELOPED-CHAR.  CHANGE OF STATE OF SKY DURING PAST HR.",
  "STATE OF SKY ON THE WHOLE UNCHANGED-CHAR. CHANGE OF THE STATE OF SKY DURING THE PAST HOUR",
  "STATE OF SKY ON THE WHOLE UNCHANGED-CHAR. CHANGE OF THE STATE OF SKY DURING THE PAST HOUR",
  "STATE OF SKY ON THE WHOLE UNCHANGED-CHAR. CHANGE OF THE STATE OF SKY DURING THE PAST HOUR",
  "CLOUDS GENERALLY FORMING OR DEVELOPING-CHAR. CHANGE OF THE STATE OF SKY DURING THE PAST HOUR",
  "RAIN",
  "STATE OF SKY ON THE WHOLE UNCHANGED-CHAR. CHANGE OF THE STATE OF SKY DURING THE PAST HOUR",
  "PRECIPITATION WITHIN SIGHT, REACHING THE GROUND OR THE SURFACE OF THE SEA, BUT DISTANT(I.E.  ESTIMATED TO BE MORE THAN 5 KM) FROM THE STATION",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "" ;

 Cloud_Type =
  "CUMULUS (CU)",
  "CUMULUS (CU)",
  "CIRRUS (CI)",
  "CUMULUS (CU)",
  "CUMULUS (CU)",
  "CUMULUS (CU)",
  "CUMULUS (CU)",
  "CUMULONIMBUS (CB)",
  "CUMULONIMBUS (CB)",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "" ;

 Cloud_Cover =
  "2 OKTAS     2/10-3/10",
  "0 (ZERO)",
  "1 OKTA OR LESS, BUT NOT ZERO    (1/10 OR LESS, BUT NOT ZERO)",
  "3 OKTAS     4/10",
  "1 OKTA OR LESS, BUT NOT ZERO    (1/10 OR LESS, BUT NOT ZERO)",
  "1 OKTA OR LESS, BUT NOT ZERO    (1/10 OR LESS, BUT NOT ZERO)",
  "1 OKTA OR LESS, BUT NOT ZERO    (1/10 OR LESS, BUT NOT ZERO)",
  "6 OKTAS     7/10-8/10",
  "1 OKTA OR LESS, BUT NOT ZERO    (1/10 OR LESS, BUT NOT ZERO)",
  "3 OKTAS     4/10",
  "3 OKTAS     4/10",
  "2 OKTAS     2/10-3/10",
  "0 (ZERO)",
  "0 (ZERO)",
  "0 (ZERO)",
  "0 (ZERO)",
  "5 OKTAS     6/10",
  "6 OKTAS     7/10-8/10",
  "8 OKTAS     10/10",
  "6 OKTAS     7/10-8/10",
  "0 (ZERO)",
  "8 OKTAS     10/10",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "" ;

 dataset =
  "bottle/rossette/net",
  "bottle/rossette/net",
  "bottle/rossette/net",
  "bottle/rossette/net",
  "bottle/rossette/net",
  "bottle/rossette/net",
  "bottle/rossette/net",
  "bottle/rossette/net",
  "bottle/rossette/net",
  "bottle/rossette/net",
  "bottle/rossette/net",
  "bottle/rossette/net",
  "bottle/rossette/net",
  "bottle/rossette/net",
  "bottle/rossette/net",
  "bottle/rossette/net",
  "bottle/rossette/net",
  "bottle/rossette/net",
  "bottle/rossette/net",
  "bottle/rossette/net",
  "bottle/rossette/net",
  "bottle/rossette/net",
  "bottle/rossette/net",
  "bottle/rossette/net",
  "bottle/rossette/net",
  "bottle/rossette/net",
  "bottle/rossette/net",
  "bottle/rossette/net",
  "bottle/rossette/net",
  "bottle/rossette/net",
  "bottle/rossette/net",
  "bottle/rossette/net",
  "bottle/rossette/net",
  "bottle/rossette/net",
  "bottle/rossette/net",
  "bottle/rossette/net",
  "bottle/rossette/net",
  "bottle/rossette/net",
  "bottle/rossette/net",
  "bottle/rossette/net",
  "bottle/rossette/net",
  "bottle/rossette/net",
  "bottle/rossette/net",
  "bottle/rossette/net",
  "bottle/rossette/net",
  "bottle/rossette/net",
  "bottle/rossette/net",
  "bottle/rossette/net",
  "bottle/rossette/net",
  "bottle/rossette/net",
  "bottle/rossette/net",
  "bottle/rossette/net",
  "bottle/rossette/net",
  "bottle/rossette/net",
  "bottle/rossette/net",
  "bottle/rossette/net",
  "bottle/rossette/net",
  "bottle/rossette/net",
  "bottle/rossette/net",
  "bottle/rossette/net",
  "bottle/rossette/net",
  "bottle/rossette/net",
  "bottle/rossette/net",
  "bottle/rossette/net",
  "bottle/rossette/net",
  "bottle/rossette/net",
  "bottle/rossette/net",
  "bottle/rossette/net",
  "bottle/rossette/net",
  "bottle/rossette/net",
  "bottle/rossette/net",
  "bottle/rossette/net",
  "bottle/rossette/net",
  "bottle/rossette/net",
  "bottle/rossette/net",
  "bottle/rossette/net",
  "bottle/rossette/net",
  "bottle/rossette/net",
  "bottle/rossette/net",
  "bottle/rossette/net",
  "bottle/rossette/net",
  "bottle/rossette/net",
  "bottle/rossette/net",
  "bottle/rossette/net",
  "bottle/rossette/net",
  "bottle/rossette/net",
  "bottle/rossette/net",
  "bottle/rossette/net",
  "bottle/rossette/net",
  "bottle/rossette/net",
  "bottle/rossette/net",
  "bottle/rossette/net",
  "bottle/rossette/net",
  "bottle/rossette/net",
  "bottle/rossette/net",
  "bottle/rossette/net",
  "bottle/rossette/net",
  "bottle/rossette/net",
  "bottle/rossette/net",
  "bottle/rossette/net",
  "bottle/rossette/net",
  "bottle/rossette/net",
  "bottle/rossette/net",
  "bottle/rossette/net",
  "bottle/rossette/net",
  "bottle/rossette/net",
  "bottle/rossette/net",
  "bottle/rossette/net",
  "bottle/rossette/net",
  "bottle/rossette/net",
  "bottle/rossette/net",
  "bottle/rossette/net",
  "bottle/rossette/net",
  "bottle/rossette/net",
  "bottle/rossette/net",
  "bottle/rossette/net",
  "bottle/rossette/net",
  "bottle/rossette/net",
  "bottle/rossette/net",
  "bottle/rossette/net",
  "bottle/rossette/net",
  "bottle/rossette/net",
  "bottle/rossette/net",
  "bottle/rossette/net",
  "bottle/rossette/net",
  "bottle/rossette/net",
  "bottle/rossette/net",
  "bottle/rossette/net",
  "bottle/rossette/net",
  "bottle/rossette/net",
  "bottle/rossette/net",
  "bottle/rossette/net",
  "bottle/rossette/net",
  "bottle/rossette/net",
  "bottle/rossette/net",
  "bottle/rossette/net",
  "bottle/rossette/net",
  "bottle/rossette/net",
  "bottle/rossette/net",
  "bottle/rossette/net",
  "bottle/rossette/net",
  "bottle/rossette/net",
  "bottle/rossette/net",
  "bottle/rossette/net",
  "bottle/rossette/net",
  "bottle/rossette/net",
  "bottle/rossette/net",
  "bottle/rossette/net",
  "bottle/rossette/net",
  "bottle/rossette/net",
  "bottle/rossette/net",
  "bottle/rossette/net",
  "bottle/rossette/net",
  "bottle/rossette/net",
  "bottle/rossette/net",
  "bottle/rossette/net",
  "bottle/rossette/net",
  "bottle/rossette/net",
  "bottle/rossette/net",
  "bottle/rossette/net",
  "bottle/rossette/net",
  "bottle/rossette/net",
  "bottle/rossette/net",
  "bottle/rossette/net",
  "CTD",
  "bottle/rossette/net",
  "bottle/rossette/net",
  "bottle/rossette/net",
  "bottle/rossette/net" ;

 Ref_Type =
  "NANSEN CAST (REVERSING THERMOMETER)",
  "NANSEN CAST (REVERSING THERMOMETER)",
  "NANSEN CAST (REVERSING THERMOMETER)",
  "NANSEN CAST (REVERSING THERMOMETER)",
  "NANSEN CAST (REVERSING THERMOMETER)",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "" ;

 Visibility =
  "insufficient information",
  "insufficient information",
  "insufficient information",
  "no fix necessary",
  "no fix necessary",
  "no fix necessary",
  "insufficient information",
  "insufficient information",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "" ;

 Absol_Humidity = _, _, _, _, _, 2.9, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, 15.2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, 2.7, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 12.9, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, 11.9, 2.6, 7.4, 7.5, _, _, _, _, 7.5, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 10.9, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, 10.9, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 dbase_orig =
  "NODC archive (1992)",
  "NODC archive (1992)",
  "NODC archive (1992)",
  "GODAR Project",
  "NODC archive (1992)",
  "GODAR Project",
  "NODC archive (1992)",
  "NODC archive (1992)",
  "NODC archive (1992)",
  "GODAR Project",
  "NODC archive (1992)",
  "NODC archive (1992)",
  "NODC archive (1992)",
  "GODAR Project",
  "GODAR Project",
  "NODC archive (1992)",
  "GODAR Project",
  "GODAR Project",
  "GODAR Project",
  "GODAR Project",
  "NODC archive (1992)",
  "NODC archive (1992)",
  "NODC archive (1992)",
  "GODAR Project",
  "NODC archive (1992)",
  "NODC archive (1992)",
  "GODAR Project",
  "NODC archive (1992)",
  "NODC archive (1992)",
  "GODAR Project",
  "GODAR Project",
  "GODAR Project",
  "GODAR Project",
  "NODC archive (1992)",
  "NODC archive (1992)",
  "NODC archive (1992)",
  "GODAR Project",
  "NODC archive (1992)",
  "GODAR Project",
  "NODC archive (1992)",
  "NODC archive (1992)",
  "GODAR Project",
  "GODAR Project",
  "GODAR Project",
  "GODAR Project",
  "NODC archive (1992)",
  "NODC archive (1992)",
  "NODC archive (1992)",
  "GODAR Project",
  "GODAR Project",
  "GODAR Project",
  "GODAR Project",
  "GODAR Project",
  "GODAR Project",
  "NODC archive (1992)",
  "NODC archive (1992)",
  "GODAR Project",
  "NODC archive (1992)",
  "GODAR Project",
  "NODC archive (1992)",
  "GODAR Project",
  "NODC archive (1992)",
  "NODC archive (1992)",
  "GODAR Project",
  "NODC archive (1992)",
  "GODAR Project",
  "NODC archive (1992)",
  "NODC archive (1992)",
  "NODC archive (1992)",
  "GODAR Project",
  "GODAR Project",
  "GODAR Project",
  "NODC archive (1992)",
  "NODC archive (1992)",
  "NODC archive (1992)",
  "NODC archive (1992)",
  "GODAR Project",
  "GODAR Project",
  "NODC archive (1992)",
  "NODC archive (1992)",
  "GODAR Project",
  "NODC archive (1992)",
  "GODAR Project",
  "NODC archive (1992)",
  "GODAR Project",
  "NODC archive (1992)",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "" ;

 z = 0, 10, 20, 30, 50, 75, 100, 125, 150, 200, 250, 300, 400, 500, 600, 700, 
    800, 900, 1000, 1100, 1200, 1300, 1400, 1500, 1750, 2000 ;

 zcast_WODflag =
  0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _,
  0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _,
  0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _,
  0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _,
  0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _,
  0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _,
  0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _,
  0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _,
  0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 Temperature =
  20.4, _, _, _, 19.85, _, 19.3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _,
  27.83, 27.76, 26.6, 25.9, 25.47, 24, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _,
  3.9, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  3.05, 3.06, 3.08, 3.2, 3.24, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _,
  2.92, 2.96, 3.09, 3.09, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2.92, 3.05, 4.35, 4.74, 4.74, 4.7, 4.71, 4.66, 4.63, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _,
  16.7, 16.58, 16.55, 16.5, 15.83, 15.32, 14.78, 14.27376, 13.87, 13.41, 
    12.88, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, 0.7164688, 0.737972, 0.7207446, 0.7788591, _, 3.157495, _, 5.772188, _, 
    8.722754, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, 0.7137667, 0.7389348, 0.7215973, 0.7611144, _, 3.120401, _, 5.736207, _, 
    8.714807, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2.76, 2.79, 2.77, 2.77, 2.77, 2.83, 2.92, 3.07, 3.34, 4.3, 3.68, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _,
  7.25, 7.259927, 7.250355, 7.24745, 7.050881, 6.96, 6.936899, 6.76267, 
    6.467665, 5.765314, 5.226902, 4.680755, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _,
  3.8, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  3.01, 2.74, 3.72, 4.01, 4.39, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _,
  17.2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  26.04, 26.04, 26.04, 26.04, 25.63268, 20.02, 17.23, 14.67063, 12.7111, 
    11.44993, 10.79198, 10.2666, 9.416855, 8.749153, _, _, _, 5.274754, 
    5.031479, 4.83399, 4.785833, _, 4.39425, _, _, _,
  14.3, 14.19, 14.01, 13.9, 13.07, 10.66, 9.68, 9.241285, 8.91, 8.33, 7.72, 
    7.25, 6.57, 5.95, 5.31, 4.825559, 4.47, 4.221797, 3.97, 3.705, 3.43, _, 
    _, _, _, _,
  3.5, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  3.5, 14.19, 14.01, 13.9, 13.07, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _,
  18.42, 18.17, 17.55, 17.34, 17.09, 16.97, 16.66, 16.60569, 16.55, 16.41, 
    15.54874, 15.10027, 13.95, 12.75, 10.87, 9.366593, 8.22, 7.5344, 
    6.978853, 6.44021, 5.95, 5.48175, 5.076794, 4.72, _, 3.9,
  17, 16.7725, 16.59947, 16.22422, 15.62345, 14.63129, 13.81432, 13.65265, 
    13.17818, _, 10.89364, 9.896256, 8.293365, _, _, _, _, _, _, _, _, _, _, 
    _, _, _,
  2.73, 2.74, 2.74, 2.74, 2.76, 2.95, 4.39, 4.42, 4.32, 3.75, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _,
  0.8, 0.7388462, 0.6776923, 0.6165385, 0.4942308, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _,
  4.4, 4.44, 4.55, 4.45, 4.37, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _,
  19.44, 19.41653, 19.41, 19.37877, 19.28085, 19.17673, 19.06, 18.74782, 
    18.5354, 17.70466, 16.89619, 16.08079, 14.14384, 11.68, 8.763053, 
    6.488856, _, 4.519095, 3.982477, 3.594397, 3.201619, 2.824135, _, _, _, _,
  27.52, 27.53, 27.52228, 27.522, 27.53, 27.47, 26.68937, 23.8807, 18.4668, 
    14.93976, 12.66838, 11.46792, 10.14188, 7.831767, 6.61, _, _, _, _, _, _, 
    _, _, _, _, _,
  3.5, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  2.55, 2.26, 3.49, 3.54, 3.88, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _,
  25.28, 24.81, 24.5166, 24.33872, 24.04076, 23.91516, 23.38256, 22.06804, 
    20.50591, 18.98648, 17.44844, 16.06879, 13.1077, 10.2208, 7.849243, _, _, 
    4.220284, 3.659655, _, 3.056614, _, _, 2.620602, _, _,
  2.66, 2.73, 3.56, 4.01, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _,
  2.41, 2.52, 2.58, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _,
  16.3, 16.07, 15.97, 15.93, 15.88, 15.4605, 14.83, 14.17349, 13.43, 12.87, 
    11.48333, 9.27, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  17, 16.82, 16.48, 16.22, 15.88, 14.99, 14.19, 13.79952, 13.34, 12.06, 
    10.85667, 9.73, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  17, 16.82, 16.48, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _,
  2.01, 2.26, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _,
  16.5, 16.24, 16.15, 16.1, 16.05, 15.76172, 15.27, 14.7841, 14.15, 12.36, 
    10.95173, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  15.35, 15.34377, 15.34, 15.34, 15.31812, 14.33694, 12.64815, 11.08958, 
    9.954114, 8.785531, 8.163257, 7.656954, 5.869786, 5.203469, _, _, _, 
    3.855511, 3.595377, 3.345377, _, _, _, _, _, _,
  5.36, 5.34, 5.34, 5.34, 5.32, 5.36, 5.39, 5.36047, 5.34, 5.36, 5.37, 5.33, 
    5.04, 4.82, 4.5, 4.18, 4.02, 3.89, 3.76, 3.629999, 3.5, 3.52353, 3.55031, 
    3.56, _, 3.320903,
  2.7, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  20.3, _, _, _, 19.6, _, 18.9, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _,
  30.17, 28.2, 26.77, 26.45481, 26.27, 26.27, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _,
  0.2, 1.2, 2.55, 5.48, 6.23, 6.46, 6.41, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _,
  0.8, _, 0.9356923, 1.003538, 1.139231, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  5.24, 5.27, 5.26, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _,
  5.23, 5.25, 5.23, 5.24, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _,
  0.3, 1.06, 1.945645, 3.603647, 6.02, 6.24, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _,
  2.2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  26.2, 26.20841, 26.22, 26.23373, 26.17361, 22.63, 15.81303, 13.35638, 
    12.60369, _, 10.82407, _, _, 7.818521, 6.869727, _, _, 5.08116, 4.948574, 
    4.826803, _, _, _, _, _, _,
  27.98, 27.98, 27.99677, 27.99731, 27.98794, 27.9148, 27.70919, 22.6878, 
    18.60445, 14.10852, 12.28513, 11.82, 10.30208, 8.361901, 7.13, _, _, _, 
    _, _, _, _, _, _, _, _,
  14.94, 14.84, 14.74, 13.94, 12.25, 11.24, 10.16, 9.647418, 9.31, 8.76, 
    8.36, 7.78, 6.97, 6.08, 5.22, 4.956587, 4.67, 4.299918, 3.92, 3.635, 
    3.41, _, _, _, _, _,
  5.27, 5.33, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _,
  2.45, 2.39, 2.46, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _,
  4.99, 5.02, 5.01, 5, 4.93, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _,
  2.56, 2.38, 3.61, 3.95, 4.04, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _,
  2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2.38, 3.61, 3.95, 4.04, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _,
  2.75, 2.75, 2.75, 2.75, 2.75, 2.94, 2.94, 2.92, 3.95, 4.42, 4.11, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _,
  25.67, 25.05762, 24.89336, 24.76658, 24.4787, 24.02281, 23.35505, 22.51032, 
    21.64579, 19.91469, 18.19936, 16.93218, 14.55191, 11.56844, _, _, _, 
    4.225826, 3.852011, 3.433742, 3.127324, _, 2.704762, _, _, _,
  0.15, 2.88, 4.52, 5.07, 6.42, 4.8, 5.56, 5.63, 5.7, 5.97, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _,
  0.15, 2.88, 4.52, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _,
  5.37, 5.47, 5.6, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _,
  5.36, 5.43, 5.66, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _,
  18, 18.02463, 18.06365, 18.10813, 18.07633, 18.06488, 17.93806, 17.58196, 
    17.3531, 17.21692, _, _, _, 12.33248, 9.497299, _, _, _, 3.991845, _, _, 
    2.918632, _, _, _, _,
  6.5, 6.240008, 6.249479, 6.241696, 6.233809, 6.245715, 6.25, 6.238973, 
    6.120853, 5.914982, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 2.846666, 4.99, 6.18, 5.97, 6.46, 5.87, 6.2, 6.61, 6.36, 6.01, 5.85, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _,
  0.9, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  2.5, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  27.91, 24.32, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _,
  22.34, 22.31837, 22.31252, 22.32657, 21.15783, 17.03691, _, _, _, _, 
    12.27514, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  5.76, 5.77, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _,
  6.58, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  0.2, 0.841114, 3.64491, 5.41, 6.53, 6.29, 6.46, 6.41, 6.26, 6.11, 5.79, 
    5.55, 5.04, _, _, _, _, _, _, _, _, _, _, _, _, _,
  5.83, 5.88, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _,
  2.6, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  15.59, 15.5409, 15.53011, 15.55197, 15.68771, 15.66187, 13.98757, 12.2025, 
    10.74217, 9.073494, 8.46131, 7.637049, 6.037966, _, _, _, _, 3.744935, 
    3.527421, _, _, _, _, _, _, _,
  1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  5.47, 5.49, 5.37, 5.26, 5.37, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _,
  5.36, 5.41, 5.46, 5.46, 5.41, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _,
  28.08, 27.86, 27.28, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _,
  2.35, 2.45, 4.35, 4.27, 3.89, 4.1, 5.04, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _,
  2.35, 2.45, 4.35, 4.27, 3.89, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _,
  2.35, 2.45, 4.35, 4.27, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _,
  6.47, 6.48, 6.49, 6.48, 6.47, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _,
  19.6, _, _, _, 18.8, _, 18, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _,
  1.7, 2.17, 4.51, 5.23, 5.98, 6.41, 6.89, 6.91, 6.53, 6.18, 5.98, 5.68, 
    5.24, 4.99, 4.91, _, _, _, _, _, _, _, _, _, _, _,
  24.84, 24.84, 24.83894, 24.82, 24.71562, 18.05014, 15.55022, 14.1662, 
    13.20238, 11.79805, 11.25666, 10.53242, 9.837049, _, _, _, _, _, _, _, _, 
    _, _, _, _, _,
  4.66, 4.64, 4.64, 4.64, 4.65, 4.66, 4.68, 4.669431, 4.66, 4.65, 4.49, 4.15, 
    4.08, 3.88, 3.9, 3.78, 3.74, 3.7, 3.66, 3.571027, 3.46, 3.474166, 
    3.495371, 3.5, _, 3.293035,
  14.48, 14.48, 14.31, 14.25, 13.8, 12.3, 10.58, 9.693413, 9.35, 9.02, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  22.06, 22.06, 22.05658, 22.05108, 22.04327, 19.43, 15.73, 14.06087, 
    13.43699, 12.65478, 11.87931, 11.59596, 10.57941, 9.776645, _, _, _, _, 
    _, _, _, _, _, _, _, _,
  17.3, 17.14, 16.99, 16.62, 13.42, 11.56, 10.68, 9.777302, 8.86, 7.52, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2.75, 2.93, 3.54, 4.28, 4.34, 4.71, 5.94, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _,
  6.6, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  2.5, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  18.96, 18.96, 18.96, 18.98737, 18.9424, 18.95927, 18.82436, 18.70539, 
    18.59475, 17.77199, 17.32032, 16.35955, 14.8558, 13.94198, 11.3478, 
    8.58965, _, 5.299035, _, 3.656482, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  7.3, 6.7, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  7.2, 6.68, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _,
  2.63, 2.63, 2.64, 2.61, 2.59, 2.59, 2.59, 3.24, 4.04, 4.11, 3.97, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _,
  2.45, 2.87, 5.28, 6.12, 5.47, 5.93, 6.48, 6.07, 6.38, 5.7, 5.94, 5.54, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _,
  6.81, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  25.44, 25.33, 25.09505, 25.04403, 24.95808, 24.89181, 24.69283, 24.51, 
    24.36559, 22.37936, 19.33206, 17.45809, 15.17424, 11.86519, 8.789974, _, 
    _, 4.480542, 3.962507, 3.526095, 3.236801, _, _, _, _, _,
  7.3, 7.03, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _,
  1.72, 2.08, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _,
  2.81, 2.81, 2.81, 2.81, 2.82, 2.86, 2.71, 2.64, 3.17, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _,
  6.81, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  26.68, 26.65783, 26.62935, 26.61464, 26.57897, 26, 20.10464, 16.31124, 
    14.41121, 11.55575, 10.65693, 9.85543, 8.628658, 7.618165, 6.807902, _, 
    _, 5.001948, 4.878128, 4.776842, 4.77, _, 4.419187, _, _, _,
  28.14, 27.98, 27.29, 25.18, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _,
  2.5, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  2.5, 27.98, 27.29, 25.18, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _,
  17.24, 17.15, 16.8, 16.67561, 16.65, 16.46, 16.2, 16.02009, 15.83, 15.41, 
    15.28677, 15.28, 14.01, 12.54, 11.24, 9.743163, 8.06, 7.588541, 7.112982, 
    6.553833, 5.99, 5.437455, 4.880647, _, _, 3.7,
  3.88, 3.82, 3.73, 3.68, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _,
  15.4, 15.35237, 15.33207, 15.33205, 15.39818, 15.45313, 13.92242, 12.33165, 
    10.75306, 8.761237, 8.121367, 7.332345, 5.814312, 4.99534, _, _, _, 
    3.826821, 3.568124, 3.366719, _, _, _, _, _, _,
  3, 2.92, 5.24, 4.71, 4.96, 4.74, 4.7, 4.7, 4.71, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _,
  0.5, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  6.93, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  6.93, 2.92, 5.24, 4.71, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _,
  27.91, 27.92, 27.41, 24.92, 23.96, 23.34, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _,
  2.44, 2.43, 2.44, 2.46, 2.44, 2.4, 2.24, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _,
  2.95, 2.61, 3.39, 5.01, 4.69, 4.55, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _,
  0.6, 0.5095745, 0.419149, 0.3287234, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _,
  19, _, _, _, 18.4, _, 17.8, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _,
  4.07, 4.007621, 3.804544, 3.71, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _,
  17.88, 17.3, 16.47, 16.22, 13.35, 11.06, 10.16, 9.378039, 8.72, 7.79, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  17.46, 17.44, 17.44, 17.47744, 17.45169, 17.47818, 17.47315, 17.3753, 
    17.35873, 17.24541, 17.13066, 16.77057, 14.86571, 12.52032, _, _, 
    5.421472, 4.618513, _, _, _, _, _, _, _, _,
  14, 14.2, 14.02, 14, 13.69, 13.03, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _,
  3.4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  3.4, 14.2, 14.02, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _,
  2.56, 2.6, 2.36, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _,
  2.85, 2.76, 2.98, 3.86, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _,
  7.15, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  6.92, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  21.54, 21.63, 21.44, 20.16, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _,
  3.2, 2.894651, 2.589302, 2.283953, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _,
  25.45, 25.45, 25.27052, 25.1625, 25.03133, 24.91178, 24.80051, 24.53319, 
    23.94676, 21.76394, 19.43494, 17.43725, 15.09128, 11.83682, 8.721209, _, 
    _, 4.443428, 4.018601, 3.620449, 3.291281, _, 2.795374, _, _, _,
  27.72, 27.71, 27.12, 25.51, 23.78, 22.62, 20.99, 19.50063, 17.85926, 16.4, 
    15.7, 14.14, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2.1, 2.13, 2.59, 2.58, 3.79, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _,
  15.58, 15.482, 15.44, 15.48971, 15.65, 15.4844, 13.41086, 11.48292, 
    9.965707, 8.590878, 8.097981, 7.501308, 6.134176, 5.529526, _, _, _, 
    3.866576, 3.617763, 3.380562, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  14.08, 14.08, 14.08, 13.98, 13.94, 13.78, 13.22, 11.35881, 9.36, 8.8, 8.08, 
    7.42, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2.2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  3.15, 3.13, 2.68, 2.95, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _,
  2.5, _, 2.468308, 2.452461, 2.420769, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _,
  28.23, 28.23, 27.18, 26.0176, 24.33, 23.07, 21.75, 19.68174, 18.62, 16.37, 
    14.82, 12.97, 11.14, 9.85, 8.07, _, _, _, _, _, _, _, _, _, _, _,
  3.6, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  3.6, 28.23, 27.18, 26.0176, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _,
  17.55, 17.5465, 17.57399, 17.55053, 17.56863, 17.55105, 17.314, 17.264, 
    17.214, 17.13718, 17.09484, 16.9427, 15.36974, 12.86661, 10.31372, _, _, 
    4.123011, 4.037994, _, 3.189087, _, _, _, _, _,
  3.4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  3.7, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  3.7, 17.5465, 17.57399, 17.55053, 17.56863, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _,
  19.4, _, _, _, 18.9, _, 18.4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _,
  2.6, _, _, _, 2.793452, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _,
  10.61, 10.60814, 10.58178, 10.59157, 10.6, 10.59787, 10.56518, 10.51874, 
    9.810402, 5.913959, 2.035888, 0.9324624, 0.4477943, 0.301725, 0.2033058, 
    _, _, _, _, _, _, _, _, _, _, _,
  13.9, 13.88247, 13.77175, 13.69722, 13.06908, 10.43856, 9.424856, 9.218444, 
    9.005425, 8.593699, 7.914983, 7.471694, 6.700624, 5.938673, _, _, _, 
    4.113402, 3.841489, 3.59319, _, _, _, _, _, _,
  3.09, 3.15, 3.54, 4.02, 4.15605, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _,
  1.34, 1.33, 1.33, 1.34, 1.35, 1.34, 1.4, 1.41, 1.46, 1.99, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _,
  25.53, 25.55, 25.54472, 25.43946, 25.21929, 24.96003, 24.72007, 24.30267, 
    23.63914, 21.43017, 19.59442, 17.73813, 14.37492, 11.15738, _, _, _, _, 
    4.170431, _, 3.374988, 3.127001, _, _, _, _,
  6.82, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  6.33, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  23.13, 23.14, 23.14, 23.13, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _,
  6.48, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  6.48, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  6.8, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  5.87, 5.86, 5.864999, 5.868706, 5.846045, 5.83, 5.743161, 5.114305, 5.121, 
    4.787252, 4.351286, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  6.58, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  7.17, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  7.13, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  6.81, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _ ;

 Temperature_sigfigs =
  3, _, _, _, 3, _, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4, 4, 4, 4, 4, 4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4, 4, 4, 4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, 3, 3, 3, 3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4, 3, 3, 3, 3, _, 4, _, 4, _, 4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4, 3, 3, 3, 3, _, 4, _, 4, _, 4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 3, 3, _, _, _, 3, 3, 3, 3, _, 3, _, _, _,
  4, 4, 4, 4, 4, 4, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, _, _, _, _, _,
  3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 4, 4, 4, 4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 3, 3, 3, 3, 3, 3, 3, 3, 3, _, 3,
  4, 4, 4, 4, 4, 4, 4, 4, 4, _, 4, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, 3, 3, 3, 3, 3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 3, 3, _, 3, 3, 3, 3, 3, _, _, _, _,
  4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 3, 3, _, _, _, _, _, _, _, _, _, _, _,
  3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 3, _, _, 3, 3, _, 3, _, _, 3, _, _,
  3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4, 4, 4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4, 4, 4, 4, 4, 4, 4, 4, 3, 3, 3, 3, 3, 3, _, _, _, 3, 3, 3, _, _, _, _, _, _,
  3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, _, 3,
  3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, _, _, _, 3, _, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4, 4, 4, 4, 4, 4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 3, 3, 3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, _, 3, 4, 4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 3, 3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4, 4, 4, 4, 4, 4, 4, 4, 4, _, 4, _, _, 3, 3, _, _, 3, 3, 3, _, _, _, _, _, _,
  4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 3, 3, _, _, _, _, _, _, _, _, _, _, _,
  4, 4, 4, 4, 4, 4, 4, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, _, _, _, _, _,
  3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, _, _, _, 3, 3, 3, 3, _, 3, _, _, _,
  2, 3, 3, 3, 3, 3, 3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4, 4, 4, 4, 4, 4, 4, 4, 4, 4, _, _, _, 4, 3, _, _, _, 3, _, _, 3, _, _, _, _,
  3, 3, 3, 3, 3, 3, 3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4, 4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4, 4, 4, 4, 4, 4, _, _, _, _, 4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4, 4, 4, 4, 4, 4, 4, 4, 4, 3, 3, 3, 3, _, _, _, _, 3, 3, _, _, _, _, _, _, _,
  4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, 3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 4, 4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, 3, 3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, _, _, _, 3, _, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _,
  4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 3, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, _, 3,
  4, 4, 4, 4, 4, 4, 4, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 3, _, _, _, _, _, _, _, _, _, _, _, _,
  4, 4, 4, 4, 4, 4, 4, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, 3, 3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 3, _, 3, _, 3, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 3, _, _, 3, 3, 3, 3, _, _, _, _, _,
  3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, 3, 3, 3, 3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 3, 3, 3, 3, _, _, 3, 3, 3, 3, _, 3, _, _, _,
  2, 4, 4, 4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, 4, 4, 4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 3, 3, 3, 3, 3, 3, 3, 3, _, _, 3,
  3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4, 4, 4, 4, 4, 4, 4, 4, 4, 3, 3, 3, 3, 3, _, _, _, 3, 3, 3, _, _, _, _, _, _,
  3, 3, 3, 3, 3, 3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 4, 4, 4, 4, 4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, 3, 3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, 3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, _, _, _, 3, _, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4, 4, 4, 4, 4, 4, 4, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, _, _, 3, 3, _, _, _, _, _, _, _, _,
  4, 4, 4, 4, 4, 4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 4, 4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4, 4, 4, 4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4, 4, 4, 4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 3, _, _, 3, 3, 3, 3, _, 3, _, _, _,
  4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4, 4, 4, 4, 4, 4, 4, 4, 3, 3, 3, 3, 3, 3, _, _, _, 3, 3, 3, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4, 4, 4, 4, 4, 4, 4, 4, 3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4, _, 4, 4, 4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 3, 3, _, _, _, _, _, _, _, _, _, _, _,
  1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, 4, 4, 4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, _, _, 3, 3, _, 3, _, _, _, _, _,
  3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 4, 4, 4, 4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, _, _, _, 3, _, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4, _, _, _, 4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  5, 5, 5, 5, 5, 5, 5, 5, 4, 4, 4, 3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _,
  4, 4, 4, 4, 4, 4, 3, 3, 3, 3, 3, 3, 3, 3, _, _, _, 3, 3, 3, _, _, _, _, _, _,
  3, 3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, 3, 3, 3, 3, 3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, _, _, _, _, 3, _, 3, 3, _, _, _, _,
  3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4, 4, 4, 4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 Temperature_WODflag =
  0, _, _, _, 0, _, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, _, 0, _, 0, _, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, _, 0, _, 0, _, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 2, 2, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, 0, 0, 0, 0, _, 0, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, _, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, 0, 0, 0, 0, 0, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, 0, 0, _, 0, _, _, 0, _, _,
  0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, 0, 0, 0, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, 0,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, 0, _, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, _, 0, _, _, 0, 0, _, _, 0, 0, 0, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _,
  0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, 0, 0, 0, 0, _, 0, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, 0, 0, _, _, _, 0, _, _, 0, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, _, _, _, _, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, 0, 0, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, 0, _, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, 0, _, 0, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 9, _, _, 0, 0, 0, 0, _, _, _, _, _,
  0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, 0, 0, 0, 0, _, 0, _, _, _,
  0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, 0,
  0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, 0, 0, 0, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, 0, _, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, 0, 0, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 9, _, _, 0, 0, 0, 0, _, 0, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, 0, 0, 0, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 3, 9, 7, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, 0, 0, _, 0, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, 0, _, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, 0, 0, 0, _, _, _, _, _, _,
  0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, 0, _, 0, 0, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 2, 2, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 Temperature_WODprofileflag = 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 
    0, 0, 0, 8, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 Temperature_Instrument =
  "CTD: TYPE UNKNOWN",
  "CTD: TYPE UNKNOWN",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "" ;

 Salinity =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  33.263, 33.353, 33.466, 33.595, 33.702, 33.971, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _,
  32.496, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _,
  33.065, 33.065, 33.088, 33.113, 33.158, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _,
  33.065, 33.065, 33.088, 33.113, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _,
  34.415, 34.416, 34.435, 34.438, 34.461, 34.485, 34.493, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _,
  32.483, 33.501, 34.3, 34.584, 34.713, 34.779, 34.784, 34.787, 34.786, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  34.796, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _,
  32.05, 32.04581, 32.04959, 32.07681, 32.29493, _, 32.74262, _, 33.19654, _, 
    34.74675, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  32.05, 32.04531, 32.05011, 32.06667, 32.28797, _, 32.73652, _, 33.18542, _, 
    34.74072, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  34.546, 34.519, 34.548, 34.549, 34.549, 34.548, 34.595, 34.634, 34.63, 
    34.928, 34.894, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  33.97, 33.967, 33.967, 33.96696, 33.96315, 33.93877, 33.93333, 33.92719, 
    33.91087, 33.84789, 33.84887, 33.90342, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _,
  32.524, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _,
  32.87, 33.11, 34.01, 34.35, 34.63, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _,
  34.792, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _,
  36.232, 36.23504, 36.241, 36.259, 36.24509, 36.072, 35.986, 35.66021, 
    35.30505, 35.11867, 34.95878, 34.95788, 34.89747, 34.88355, _, _, _, 
    34.68987, 34.71536, 34.76029, 34.83894, _, 34.91093, _, _, _,
  33.07, 33.13, 33.13, 33.13, 33.22, 33.38, 33.59, 33.73714, 33.83, 33.95, 
    34.01, 34.03, 34.11, 34.14, 34.2, 34.25075, 34.29, 34.30759, 34.33, 
    34.35751, 34.39, _, _, _, _, _,
  32.34, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  32.34, 33.13, 33.13, 33.13, 33.22, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _,
  36.402, 36.382, 36.378, 36.37, 36.37, 36.358, 36.32, 36.30083, 36.298, 
    36.332, 35.97274, 36.08452, 35.926, 35.749, 35.502, 35.35541, 35.295, 
    35.34646, 35.38752, 35.33565, 35.27, 35.21878, 35.17654, 35.143, _, 35.072,
  34.776, 34.74215, 34.76275, 34.76781, 34.73405, 34.66456, 34.60972, 
    34.58268, 34.55399, _, 34.43925, 34.3874, 34.31, _, _, _, _, _, _, _, _, 
    _, _, _, _, _,
  34.486, 34.492, 34.486, 34.487, 34.488, 34.601, 34.792, 34.871, 34.938, 
    34.903, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  31.47, 31.56731, 31.66462, 31.76192, 31.95654, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _,
  33.325, 33.333, 33.327, 33.338, 33.329, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _,
  34.819, 34.818, 34.8186, 34.81957, 34.8224, 34.824, 34.824, 34.82389, 
    34.82281, 34.75211, 34.71763, 34.67879, 34.5493, 34.351, 34.15464, 
    34.21729, _, 34.22391, 34.24609, 34.30987, 34.37477, 34.45275, _, _, _, _,
  35.4, 35.4, 35.38534, 35.38, 35.38, 35.4, 35.52759, 35.51575, 35.27435, 
    35.09121, 34.90088, 34.82701, 34.75795, 34.62385, 34.57, _, _, _, _, _, 
    _, _, _, _, _, _,
  32.335, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _,
  32.85, 32.89, 34.08, 34.17, 34.33, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _,
  35.045, 35.039, 35.01566, 34.98843, 34.98246, 34.97676, 34.93372, 34.94043, 
    34.96147, 34.89981, 34.77997, 34.69369, 34.48445, 34.28025, 34.19364, _, 
    _, 34.34784, 34.40983, _, 34.50235, _, _, 34.57471, _, _,
  32.73, 33.11, 33.9, 34.28, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _,
  32.287, 33.097, 33.128, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _,
  34.788, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _,
  34.764, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _,
  34.764, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _,
  33.16, 33.26, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _,
  34.768, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _,
  33.339, 33.33739, 33.3372, 33.33742, 33.34486, 33.41191, 33.4111, 33.41358, 
    33.43826, 33.68825, 33.97136, 34.00964, 34.00618, 34.08403, _, _, _, 
    34.40784, 34.44603, 34.47663, _, _, _, _, _, _,
  34.93, 34.93, 34.92, 34.92, 34.92, 34.93, 34.92, 34.92, 34.92, 34.93, 
    34.93, 34.93, 34.91, 34.92, 34.93, 34.92, 34.93, 34.928, 34.92, 34.91066, 
    34.9, 34.916, 34.93591, 34.95, _, 34.95998,
  31.93, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  31.93, 34.93, 34.92, 34.92, 34.92, 34.93, 34.92, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _,
  32.761, 33.167, 33.552, 33.59095, 33.62881, 33.643, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _,
  22.51, 28.87, 30.61, 33.64, 34.21, 34.36, 34.39, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _,
  31.284, _, 31.57415, 31.71923, 32.00938, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _,
  34.41, 34.419, 34.472, 34.461, 34.475, 34.49, 34.504, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _,
  34.852, 34.858, 34.879, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _,
  34.855, 34.861, 34.878, 34.86, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _,
  25.86, 29.19, 30.58, 33.61, 34.21, 34.48, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _,
  31.788, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _,
  36.148, 36.1445, 36.141, 36.15512, 36.17776, 36.183, 35.83249, 35.52404, 
    35.30489, _, 35.02707, _, _, 34.7343, 34.66538, _, _, 34.6242, 34.68884, 
    34.75538, _, _, _, _, _, _,
  35.51, 35.51, 35.51, 35.51, 35.51045, 35.53, 35.53857, 35.64729, 35.40662, 
    35.0468, 34.88926, 34.86, 34.80188, 34.66204, 34.6, _, _, _, _, _, _, _, 
    _, _, _, _,
  33.13, 33.14, 33.13, 33.15, 33.31, 33.38, 33.52, 33.61072, 33.69, 33.84, 
    33.93, 33.96, 34.01, 34.05, 34.06, 34.1737, 34.28, 34.3041, 34.33, 
    34.3625, 34.4, _, _, _, _, _,
  34.83, 34.89, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _,
  33.091, 33.091, 33.172, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _,
  33.508, 33.515, 33.505, 33.507, 33.549, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _,
  32.785, 32.834, 34.145, 34.325, 34.377, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _,
  31.795, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _,
  31.795, 32.834, 34.145, 34.325, 34.377, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _,
  34.331, 34.332, 34.33, 34.332, 34.337, 34.413, 34.487, 34.524, 34.649, 
    34.852, 34.912, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  34.921, 34.94062, 34.92959, 34.93235, 34.933, 34.93653, 34.937, 34.937, 
    34.937, 34.91289, 34.81304, 34.73428, 34.56062, 34.34695, _, _, _, 
    34.33322, 34.40514, 34.45682, 34.49522, _, 34.55121, _, _, _,
  25.65, 31.55, 33.39, 33.95, 34.44, 34.418, 34.62, 34.687, 34.71, 34.78, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  25.65, 31.55, 33.39, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _,
  34.89, 34.9, 34.93, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _,
  34.89, 34.92, 34.96, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _,
  34.868, 34.83327, 34.835, 34.835, 34.84614, 34.83987, 34.81302, 34.8237, 
    34.83521, 34.84086, _, _, _, 34.52201, 34.31454, _, _, _, 34.29376, _, _, 
    34.40644, _, _, _, _,
  35.186, 35.17584, 35.16713, 35.15984, 35.14954, 35.146, 35.1471, 35.1505, 
    35.15607, 35.15713, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  24.55, 31.21, 33.8, 34.3, 34.47, 34.73, 34.74, 34.866, 34.99, 35.02, 
    35.032, 35.028, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  31.512, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _,
  31.868, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _,
  33.82, 35.17, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _,
  35.62, 35.62, 35.62201, 35.65499, 35.66625, 35.58521, _, _, _, _, 35.01934, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  34.94, 34.95, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _,
  33.95, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  25.28, 26.74, 33.79, 34.29, 34.73, 34.827, 34.92, 34.982, 34.98, 35.02, 
    35.014, 35.006, 34.98, _, _, _, _, _, _, _, _, _, _, _, _, _,
  34.97, 35, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _,
  32.039, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _,
  33.54, 33.5371, 33.53774, 33.53844, 33.58583, 33.65594, 33.65178, 33.63589, 
    33.62712, 33.77096, 33.95632, 33.98427, 33.947, _, _, _, _, 34.37587, 
    34.43224, _, _, _, _, _, _, _,
  31.897, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _,
  33.843, 33.848, 33.867, 33.875, 33.901, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _,
  33.65, 33.66536, 33.6965, 33.718, 33.858, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _,
  35.19, 35.19, 35.23, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _,
  32.05, 32.74, 34.38, 34.43, 34.45, 34.51, 34.74, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _,
  32.05, 32.74, 34.38, 34.43, 34.45, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _,
  32.05, 32.74, 34.38, 34.43, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _,
  35.11, 35.15, 35.139, 35.128, 35.142, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _,
  35.11, 35.15, 35.139, 35.128, 35.142, 34.51, 34.74, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _,
  29.15, 30.63, 33.08, 33.86, 34.32, 34.65, 34.88, 34.976, 34.99, 35.01, 
    35.006, 35.002, 34.98, 34.966, 34.96, _, _, _, _, _, _, _, _, _, _, _,
  35.97, 36.03, 36, 36, 36, 35.98263, 35.74224, 35.51525, 35.33751, 35.17077, 
    35.13744, 35.01161, 34.99259, _, _, _, _, _, _, _, _, _, _, _, _, _,
  34.87, 34.87, 34.87, 34.86, 34.86, 34.87, 34.86, 34.86616, 34.87, 34.86, 
    34.86, 34.85, 34.86, 34.86, 34.88, 34.89, 34.89, 34.89, 34.89, 34.89, 
    34.89, 34.90047, 34.91055, 34.92, _, 34.94986,
  33.05, 33.03, 33.02, 33.02, 33.16, 33.32, 33.51, 33.63588, 33.7, 33.78, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  31.839, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _,
  35.971, 35.971, 35.97076, 35.9702, 35.9734, 36.306, 35.791, 35.5155, 
    35.43669, 35.36972, 35.31249, 35.32742, 35.22511, 35.21402, _, _, _, _, 
    _, _, _, _, _, _, _, _,
  35.971, 35.971, 35.97076, 35.9702, 35.9734, 36.306, 35.791, 35.5155, 
    35.43669, 35.36972, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  32.5, 33.58, 33.94, 34.25, 34.43, 34.53, 34.853, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _,
  33.88, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  32.147, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _,
  34.837, 34.826, 34.822, 34.82053, 34.8418, 34.82808, 34.83064, 34.85067, 
    34.8325, 34.77962, 34.77356, 34.70612, 34.57946, 34.51525, 34.37948, 
    34.18861, _, 34.12378, _, 34.19843, _, _, _, _, _, _,
  34.435, 34.448, 34.459, 34.467, 34.473, 34.482, 34.505, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _,
  12.27, 12.4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _,
  12.4, 12.52, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _,
  34.378, 34.372, 34.377, 34.437, 34.447, 34.449, 34.451, 34.596, 34.72, 
    34.881, 34.873, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  30.97, 32.03, 33.85, 34.24, 34.41, 34.7, 34.93, 34.919, 34.98, 34.9, 
    35.026, 35.006, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  34.3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  34.921, 34.925, 34.97651, 34.97264, 34.96805, 34.97095, 34.96884, 34.96121, 
    34.94664, 35.01228, 34.87659, 34.7562, 34.61486, 34.36679, 34.19606, _, 
    _, 34.31483, 34.38914, 34.44161, 34.48131, _, _, _, _, _,
  12.4, 12.52, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _,
  25.592, 32.511, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _,
  34.304, 34.298, 34.302, 34.301, 34.303, 34.399, 34.426, 34.451, 34.548, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  34.09, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  36.096, 36.11409, 36.10468, 36.11569, 36.10202, 36.108, 36.15451, 35.83659, 
    35.53541, 35.18436, 34.99174, 34.95092, 34.84904, 34.77341, 34.70456, _, 
    _, 34.703, 34.703, 34.77979, 34.924, _, 34.985, _, _, _,
  35.2, 35.18, 35.21, 35.32, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _,
  32.081, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _,
  32.081, 35.18, 35.21, 35.32, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _,
  36.257, 36.254, 36.225, 36.215, 36.25, 36.239, 36.244, 36.21608, 36.177, 
    36.091, 36.05392, 36.059, 35.845, 35.658, 35.496, 35.34467, 35.221, 
    35.25654, 35.25962, 35.25241, 35.214, 35.15439, 35.06834, _, _, 34.936,
  33.398, 33.395, 33.394, 33.418, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _,
  33.389, 33.38963, 33.39, 33.39, 33.40155, 33.612, 33.49345, 33.55778, 
    33.6205, 33.76773, 33.96255, 33.97982, 33.98566, 34.04355, _, _, _, 
    34.38891, 34.43211, 34.46798, _, _, _, _, _, _,
  31.97, 33.04, 33.99, 34.31, 34.61, 34.663, 34.74, 34.744, 34.75, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  31.643, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _,
  34.22, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  34.22, 33.04, 33.99, 34.31, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _,
  35.19, 35.2, 35.2, 35.27, 35.36, 35.36, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _,
  34.278, 34.271, 34.281, 34.278, 34.281, 34.259, 34.275, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _,
  32.96, 33.2, 33.7, 34.42, 34.61, 34.65, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _,
  31.215, 31.26351, 31.31202, 31.36053, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _,
  31.215, 31.26351, 31.31202, 31.36053, 34.61, 34.65, 34.275, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  33.408, 33.39677, 33.39, 33.419, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _,
  33.408, 33.39677, 33.39, 33.419, 34.61, 34.65, 34.275, 34.744, 34.75, 
    33.76773, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  34.773, 34.773, 34.773, 34.77489, 34.77243, 34.7687, 34.77403, 34.77085, 
    34.76637, 34.76431, 34.75669, 34.70753, 34.55811, 34.39391, _, _, 
    34.06273, 34.12361, 34.20846, 34.33813, _, 34.39328, _, _, _, _,
  32.51, 33.05, 33.17, 33.18, 33.21, 33.36, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _,
  32.146, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _,
  32.146, 33.05, 33.17, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _,
  32.9, 32.894, 33.085, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _,
  32.8, 32.93, 33.33, 34.08, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _,
  34.44, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  34.2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  36.19, 36.345, 36.317, 36.388, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _,
  31.722, 31.77223, 31.82247, 31.8727, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _,
  34.968, 34.9661, 34.966, 34.96758, 34.968, 34.96929, 34.97247, 34.9767, 
    34.98168, 34.9691, 34.87401, 34.75906, 34.59373, 34.38068, 34.2073, _, _, 
    34.32797, 34.39006, 34.44788, 34.48594, _, 34.53988, _, _, _,
  35.15, 35.14, 35.18, 35.29, 35.36, 35.37, 35.38, 35.33228, 35.34776, 35.32, 
    35.3, 35.22, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  33.18, 33.17, 33.44, 33.56, 34.23, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _,
  33.363, 33.3635, 33.364, 33.42676, 33.542, 33.65202, 33.53774, 33.4374, 
    33.37753, 33.7355, 33.94806, 34.00103, 34.00443, 34.09719, _, _, _, 
    34.36185, 34.41535, 34.45923, _, _, _, _, _, _,
  34.435, 34.434, 34.433, 34.433, 34.438, 34.404, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _,
  32.75, 33.17, 33.18, 33.19, 33.2, 33.26, 33.34, 33.54372, 33.74, 33.93, 
    34.05, 34.09, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  32.415, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _,
  33.029, 33.025, 33.009, 33.151, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _,
  31.904, _, 31.95262, 31.97692, 32.02554, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _,
  35.17, 35.17, 35.16, 35.26952, 35.34, 35.34, 35.39, 35.38, 35.48, 35.45, 
    35.36, 35.14, 34.98, 34.84, 34.71, _, _, _, _, _, _, _, _, _, _, _,
  32.442, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _,
  32.442, 35.17, 35.16, 35.26952, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _,
  34.781, 34.77781, 34.776, 34.776, 34.776, 34.77335, 34.7684, 34.765, 
    34.765, 34.76489, 34.75927, 34.74256, 34.61111, 34.43912, 34.29678, _, _, 
    34.03275, 34.16891, _, 34.29655, _, _, _, _, _,
  32.39, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  32.554, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _,
  32.554, 34.77781, 34.776, 34.776, 34.776, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _,
  32.554, 34.77781, 34.776, 34.776, 34.776, 34.77335, 34.7684, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  31.942, _, _, _, 32.14914, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _,
  34.46, 34.4581, 34.43277, 34.45, 34.4507, 34.46, 34.45933, 34.45242, 
    34.40278, 34.20961, 34.10746, 34.08065, 34.0985, 34.10818, 34.11727, _, 
    _, _, _, _, _, _, _, _, _, _,
  33.2, 33.17041, 33.18105, 33.19547, 33.30012, 33.49266, 33.58032, 33.75546, 
    33.88271, 33.99828, 34.07689, 34.09967, 34.15783, 34.19337, _, _, _, 
    34.41063, 34.45155, 34.45485, _, _, _, _, _, _,
  32.268, 32.55, 32.942, 33.313, 33.39757, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _,
  34.185, 34.184, 34.184, 34.185, 34.185, 34.183, 34.187, 34.197, 34.204, 
    34.351, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  34.933, 34.933, 34.93366, 34.9453, 34.97375, 34.96835, 34.94356, 34.91057, 
    34.87083, 34.88771, 34.86363, 34.74773, 34.51406, 34.30439, _, _, _, _, 
    34.41173, _, 34.48483, 34.49783, _, _, _, _,
  35.04, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  34.31, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  35.993, 36.043, 35.986, 35.987, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _,
  34.68, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  34.68, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  35.05, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  32.62, 32.62, 32.62, 32.62, 32.62, 32.62, 32.75245, 33.48049, 33.704, 
    33.82085, 33.87206, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  34.89, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  35.05, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  35.13, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  35.1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _ ;

 Salinity_sigfigs =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  5, 5, 5, 5, 5, 5, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  5, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  5, 5, 5, 5, 5, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  5, 5, 5, 5, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  5, 5, 5, 5, 5, 5, 5, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  5, 5, 5, 5, 5, 5, 5, 5, 5, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  5, 5, 5, 5, 5, _, 5, _, 5, _, 5, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  5, 5, 5, 5, 5, _, 5, _, 5, _, 5, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  5, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  5, 5, 5, 5, 5, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  5, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, _, _, _, 5, 5, 5, 5, _, 5, _, _, _,
  4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, _, _, _, _, _,
  4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4, 4, 4, 4, 4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, _, 5,
  5, 5, 5, 5, 5, 5, 5, 5, 5, _, 5, 5, 5, _, _, _, _, _, _, _, _, _, _, _, _, _,
  5, 5, 5, 5, 5, 5, 5, 5, 5, 5, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  5, 5, 5, 5, 5, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  5, 5, 5, 5, 5, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, _, 5, 5, 5, 5, 5, _, _, _, _,
  4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, _, _, _, _, _, _, _, _, _, _, _,
  4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  5, 5, 5, 5, 5, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, _, _, 5, 5, _, 5, _, _, 5, _, _,
  5, 5, 5, 5, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 5, 5, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4, 4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, _, _, _, 5, 5, 5, _, _, _, _, _, _,
  4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, _, 4,
  4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4, 4, 4, 4, 4, 4, 4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  5, 5, 5, 5, 5, 5, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4, 4, 4, 4, 4, 4, 4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  5, _, 5, 5, 5, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  5, 5, 5, 5, 5, 5, 5, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  5, 5, 5, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  5, 5, 5, 5, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4, 4, 4, 4, 4, 4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  5, 5, 5, 5, 5, 5, 5, 5, 5, _, 5, _, _, 5, 5, _, _, 5, 5, 5, _, _, _, _, _, _,
  4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, _, _, _, _, _, _, _, _, _, _, _,
  4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, _, _, _, _, _,
  4, 4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 5, 5, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  5, 5, 5, 5, 5, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  5, 5, 5, 5, 5, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  5, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  5, 5, 5, 5, 5, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, _, _, _, 5, 5, 5, 5, _, 5, _, _, _,
  5, 5, 5, 5, 5, 5, 5, 5, 5, 5, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  5, 5, 5, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4, 4, 4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4, 4, 4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  5, 5, 5, 5, 5, 5, 5, 5, 5, 5, _, _, _, 5, 5, _, _, _, 5, _, _, 5, _, _, _, _,
  2, 5, 5, 5, 5, 5, 5, 5, 5, 5, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  5, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  5, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4, 4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  5, 5, 5, 5, 5, 5, _, _, _, _, 5, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4, 4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4, 4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, _, _, _, _, 5, 5, _, _, _, _, _, _, _,
  5, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 5, 5, 5, 5, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  5, 5, 5, 5, 5, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 4, 4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  5, 5, 5, 5, 5, 5, 5, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  5, 5, 5, 5, 5, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  5, 5, 5, 5, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  5, 5, 5, 5, 5, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  5, 5, 5, 5, 5, 5, 5, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, _, _, _, _, _, _, _, _, _, _, _,
  4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, _, 4,
  4, 4, 4, 4, 4, 4, 4, 4, 4, 4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  5, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, _, _, _, _, _, _, _, _, _, _, _, _,
  5, 5, 5, 5, 5, 5, 5, 5, 5, 5, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  5, 5, 5, 5, 5, 5, 5, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  5, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  5, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, _, 5, _, 5, _, _, _, _, _, _,
  5, 5, 5, 5, 5, 5, 5, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4, 4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4, 4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  5, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, _, _, 5, 5, 5, 5, _, _, _, _, _,
  4, 4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  5, 5, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  5, 5, 5, 5, 5, 5, 5, 5, 5, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  5, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, _, _, 5, 5, 5, 5, _, 5, _, _, _,
  2, 4, 4, 4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 4, 4, 4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, _, _, 5,
  5, 5, 5, 5, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, _, _, _, 5, 5, 5, _, _, _, _, _, _,
  5, 5, 5, 5, 5, 5, 5, 5, 5, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  5, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  5, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  5, 5, 5, 5, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 4, 4, 4, 4, 4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  5, 5, 5, 5, 5, 5, 5, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4, 4, 4, 4, 4, 4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  5, 5, 5, 5, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  5, 5, 5, 5, 4, 4, 5, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  5, 5, 5, 5, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  5, 5, 5, 5, 4, 4, 5, 5, 5, 5, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, _, _, 5, 5, 5, 5, _, 5, _, _, _, _,
  4, 4, 4, 4, 4, 4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4, 4, 4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  5, 5, 5, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4, 4, 4, 4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  5, 5, 5, 5, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  5, 5, 5, 5, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, _, _, 5, 5, 5, 5, _, 5, _, _, _,
  4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4, 4, 4, 4, 4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, _, _, _, 5, 5, 5, _, _, _, _, _, _,
  5, 5, 5, 5, 5, 5, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  5, 5, 5, 5, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  5, _, 5, 5, 5, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, _, _, _, _, _, _, _, _, _, _, _,
  2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 4, 4, 4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, _, _, 5, 5, _, 5, _, _, _, _, _,
  5, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  5, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  5, 5, 5, 5, 5, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  5, 5, 5, 5, 5, 5, 5, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  5, _, _, _, 5, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, _, _, _, _, _, _, _, _, _, _, _,
  4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, _, _, _, 4, 4, 4, _, _, _, _, _, _,
  5, 5, 5, 5, 5, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  5, 5, 5, 5, 5, 5, 5, 5, 5, 5, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, _, _, _, _, 5, _, 5, 5, _, _, _, _,
  5, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  5, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  5, 5, 5, 5, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  5, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  5, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  5, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  5, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  5, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  5, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  5, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 Salinity_WODflag =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, _, 0, _, 0, _, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, _, 0, _, 0, _, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 2, 2, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, 0, 0, 0, 0, _, 0, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 3, 6, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, _, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, _, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, 0, 0, 0, 0, 0, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, 0, 0, _, 0, _, _, 0, _, _,
  0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, 0, 0, 0, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, 0,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  5, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  8, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 5, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 5, 5, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, _, 0, _, _, 0, 0, _, _, 0, 0, 0, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 9, 0, 0, 3, 3, 6, _, _, _, _, _,
  5, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, 0, 0, 0, 0, _, 0, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, 0, 0, _, _, _, 0, _, _, 0, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, _, _, _, _, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, 0, 0, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 6, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, 0, _, 9, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, 0, 0, 0, 0, _, _, _, _, _,
  0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, 0, 0, 0, 0, _, 0, _, _, _,
  0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, 0,
  0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, 0, 0, 0, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, 0, 0, 0, 0, _, 0, _, _, _, _,
  0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, 0, 0, 0, 0, _, 0, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  5, 5, 5, 5, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, 0, 0, 0, _, _, _, _, _, _,
  0, 0, 0, 0, 8, 8, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, 0, 0, _, 0, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, 0, 0, 0, _, _, _, _, _, _,
  0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 3, 9, 9, 9, 9, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, 0, _, 0, 7, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 2, 2, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 Salinity_WODprofileflag = _, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 5, 0, 0, 0, 0, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 5, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0 ;

 Salinity_Instrument =
  "CTD: TYPE UNKNOWN",
  "CTD: TYPE UNKNOWN",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "" ;

 Oxygen =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  7.680319, 7.702711, 7.590753, 7.41162, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _,
  7.51, 7.8, 7.816203, 7.820605, 7.83, 7.835, 7.84, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _,
  7.51, 7.8, 7.816203, 7.820605, 7.83, 7.835, 7.84, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _,
  7.51, 7.8, 7.816203, 7.820605, 7.83, 7.835, 7.84, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _,
  7.51, 7.8, 7.816203, 7.820605, 7.83, 7.835, 7.84, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _,
  7.51, 7.8, 7.816203, 7.820605, 7.83, 7.835, 7.84, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _,
  7.51, 7.8, 7.816203, 7.820605, 7.83, 7.835, 7.84, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _,
  6.44, 6.469748, 6.46777, 6.406408, 6.307815, 6.289983, _, _, _, _, 4.84739, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  6.44, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  6.44, 6.469748, 6.46777, 6.406408, 6.307815, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _,
  6.44, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  6.44, 6.469748, 6.46777, 6.406408, 6.307815, 6.289983, _, _, _, _, 4.84739, 
    _, _, _, _, _, _, 0.5082346, 0.5989192, 0.6816325, _, _, _, _, _, _,
  5.99, 5.982666, 5.93, 5.852065, 5.5, 4.454475, 3.37, _, 2.286666, 2.25, _, 
    _, _, 0.61, _, _, 0.39, 0.4362669, 0.53, 0.6299999, 0.75, _, _, _, _, _,
  5.99, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  5.99, 5.982666, 5.93, 5.852065, 5.5, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _,
  5.52, 4.86, 5.68, 5.69, 5.55, 5.43, 5.39, 5.349999, 5.31, 4.84, _, _, _, 
    4.42, _, _, 3.99, 4.220038, 4.662897, _, _, _, _, 5.34, _, 5.81,
  5.52, 4.86, 5.68, 5.69, 5.55, 5.43, 5.39, 5.349999, 5.31, 4.84, _, _, _, 
    4.42, _, _, _, _, _, _, _, _, _, _, _, _,
  5.52, 4.86, 5.68, 5.69, 5.55, 5.43, 5.39, 5.349999, 5.31, 4.84, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _,
  5.52, 4.86, 5.68, 5.69, 5.55, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _,
  5.52, 4.86, 5.68, 5.69, 5.55, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _,
  5.31, 5.350178, 5.384214, 5.412107, 5.456058, 5.457073, 5.4, 5.327395, 
    5.245568, 4.887111, _, _, _, 4.28, _, _, _, _, 1.842134, 1.486485, _, _, 
    _, _, _, _,
  4.6, 4.59, 4.582742, 4.577362, 4.57, 4.52, 4.103745, 3.397454, 3.372374, 
    3.298655, 2.86512, 1.474111, 1.357624, 1.3025, 1.66, _, _, _, _, _, _, _, 
    _, _, _, _,
  4.6, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  4.6, 4.59, 4.582742, 4.577362, 4.57, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _,
  4.6, 4.59, 4.582742, 4.577362, 4.57, 4.52, 4.103745, 3.397454, 3.372374, 
    3.298655, 2.86512, 1.474111, 1.357624, 1.3025, 1.66, _, _, _, 1.842134, 
    1.486485, _, _, _, _, _, _,
  4.6, 4.59, 4.582742, 4.577362, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _,
  7.77, 7.64, 7.69, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _,
  7.77, 7.64, 7.69, 4.577362, 4.57, 4.52, 4.103745, 3.397454, 3.372374, 
    3.298655, 2.86512, 1.474111, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  7.77, 7.64, 7.69, 4.577362, 4.57, 4.52, 4.103745, 3.397454, 3.372374, 
    3.298655, 2.86512, 1.474111, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  7.77, 7.64, 7.69, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _,
  7.77, 7.64, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _,
  7.77, 7.64, 7.69, 4.577362, 4.57, 4.52, 4.103745, 3.397454, 3.372374, 
    3.298655, 2.86512, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  5.63, 5.621905, 5.613775, 5.605611, 5.589175, 5.568555, 5.507297, 5.102937, 
    4.699163, _, 3.964, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  6.74, 6.75, 6.59, 6.71, 6.73, 6.74, 6.71, 6.717522, 6.74, 6.61, 6.74, 6.62, 
    6.32, 5.88, 5.79, 5.99, 6.03, 6.156742, 6.27, 6.369616, 6.41, 6.323079, 
    6.145767, 6.07, _, 6.258677,
  6.74, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  6.74, 6.75, 6.59, 6.71, 6.73, 6.74, 6.71, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _,
  6.74, 6.75, 6.59, 6.71, 6.73, 6.74, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _,
  6.74, 6.75, 6.59, 6.71, 6.73, 6.74, 6.71, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _,
  6.74, 6.75, 6.59, 6.71, 6.73, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _,
  6.74, 6.75, 6.59, 6.71, 6.73, 6.74, 6.71, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _,
  6.74, 6.75, 6.59, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _,
  6.74, 6.75, 6.59, 6.71, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _,
  6.74, 6.75, 6.59, 6.71, 6.73, 6.74, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _,
  6.74, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  4.66, 4.66971, 4.79, 4.991245, 5.070158, 4.39, 3.299366, _, 3.214062, _, 
    3.360668, _, _, 2.323093, _, _, _, 3.268413, 3.373248, _, _, _, _, _, _, _,
  4.59, 4.68, 4.625697, 4.580917, 4.528395, 4.517986, 4.420619, 3.487561, 
    3.175897, 3.18259, 2.605351, 1.84, 1.76233, 1.916768, 1.32, _, _, _, _, 
    _, _, _, _, _, _, _,
  5.67, 5.75, 5.83, 5.394752, 4.58, 3.906068, 3.55, _, 2.873333, 2.55, _, _, 
    _, 0.69, _, _, 0.38, 0.4034031, 0.48, 0.59, 0.74, _, _, _, _, _,
  5.67, 5.75, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _,
  7.75, 7.71, 7.6, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _,
  7.75, 7.71, 7.6, 5.394752, 4.58, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _,
  7.75, 7.71, 7.6, 5.394752, 4.58, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _,
  7.75, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  7.75, 7.71, 7.6, 5.394752, 4.58, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _,
  7.75, 7.71, 7.6, 5.394752, 4.58, 3.906068, 3.55, _, 2.873333, 2.55, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  7.75, 7.71, 7.6, 5.394752, 4.58, 3.906068, 3.55, _, 2.873333, 2.55, _, _, 
    _, 0.69, _, _, 0.38, 0.4034031, 0.48, 0.59, 0.74, _, _, _, _, _,
  7.75, 7.71, 7.6, 5.394752, 4.58, 3.906068, 3.55, _, 2.873333, 2.55, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  7.75, 7.71, 7.6, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _,
  7.75, 7.71, 7.6, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _,
  7.75, 7.71, 7.6, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _,
  5.5, 5.464151, 5.438803, 5.423955, 5.426254, 5.518885, 5.459497, 5.312039, 
    5.24381, 5.247089, _, _, _, _, _, _, _, _, 2.010204, _, _, _, _, _, _, _,
  5.5, 5.464151, 5.438803, 5.423955, 5.426254, 5.518885, 5.459497, 5.312039, 
    5.24381, 5.247089, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, 6.11, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4.8, 3.221569, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _,
  4.8, 3.221569, _, _, _, _, _, _, _, _, _, 6.11, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _,
  4.8, 3.221569, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _,
  4.8, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  _, _, _, _, _, _, _, _, _, _, _, 6.22, 6.63, _, _, _, _, _, _, _, _, _, _, 
    _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  5.58, 5.574667, 5.568053, 5.560161, 5.541227, 5.512252, 5.444135, 5.341864, 
    5.208907, 4.840404, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  5.58, 5.574667, 5.568053, 5.560161, 5.541227, 5.512252, 5.444135, 5.341864, 
    5.208907, 4.840404, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  7.74, 7.74, 7.67, 7.63, 7.44, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _,
  7.76, 7.772115, 7.847106, 7.71, 8.08, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _,
  4.31, 4.55, 4.4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _,
  4.31, 4.55, 4.4, 7.71, 8.08, 5.512252, 5.444135, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _,
  4.31, 4.55, 4.4, 7.71, 8.08, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _,
  4.31, 4.55, 4.4, 7.71, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _,
  4.31, 4.55, 4.4, 7.71, 8.08, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _,
  4.31, 4.55, 4.4, 7.71, 8.08, 5.512252, 5.444135, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, 5.4, 6.51, 6.69, 6.75, _, _, _, _, _, _, 
    _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, 5.4, 6.51, _, _, _, _, _, _, _, _, _, _, 
    _, _, _,
  6.7, 6.79, 6.85, 6.75, 6.75, 6.8, 6.75, 6.75, 6.75, 6.76, 6.35, 6.68, 6.37, 
    6.36, 6.29, 6.25, 6.31, 6.28, 6.25, 6.309167, 6.37, 6.333988, 6.297238, 
    6.27, _, 6.308656,
  5.9, 5.92, 5.94, 5.82224, 5.38, 4.586572, 3.68, _, 3.26, 2.84, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _,
  5.9, 5.92, 5.94, 5.82224, 5.38, 4.586572, 3.68, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _,
  5.9, 5.92, 5.94, 5.82224, 5.38, 4.586572, 3.68, _, 3.26, 2.84, 6.35, 6.68, 
    6.37, 6.36, _, _, _, _, _, _, _, _, _, _, _, _,
  5.9, 5.92, 5.94, 5.82224, 5.38, 4.586572, 3.68, _, 3.26, 2.84, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _,
  5.9, 5.92, 5.94, 5.82224, 5.38, 4.586572, 3.68, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _,
  5.9, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  5.9, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  5.5, 5.46301, 5.434524, 5.414541, 5.400101, 5.446808, 5.496724, 5.413118, 
    5.235168, 4.683627, _, _, _, _, _, _, _, 3.10422, _, _, _, _, _, _, _, _,
  5.5, 5.46301, 5.434524, 5.414541, 5.400101, 5.446808, 5.496724, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  5.5, 5.46301, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _,
  5.5, 5.46301, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _,
  5.5, 5.46301, 5.434524, 5.414541, 5.400101, 5.446808, 5.496724, 5.413118, 
    5.235168, 4.683627, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, 6.27, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, 6.27, _, _, _, _, _, 3.10422, _, _, _, _, 
    _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, 6.27, _, _, _, _, _, 3.10422, _, _, _, _, 
    _, _, _, _,
  4.47, 4.7, 4.78, 4.86, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _,
  4.47, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  4.47, 4.7, 4.78, 4.86, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _,
  5.68, 6.33, 5.65, 5.5084, 5.38, 5.14, 5.24, 5.259109, 5.28, 5.34, _, 
    5.133849, 4.66, 4.52, _, _, 4.04, 4.099923, 4.306094, _, _, _, _, _, _, 
    5.98,
  7.53, 7.58, 7.51, 7.51, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _,
  5.62, 5.608697, 5.600054, 5.594069, 5.590138, 5.60521, 5.594419, 5.387138, 
    5.139074, _, 4.107687, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  5.62, 5.608697, 5.600054, 5.594069, 5.590138, 5.60521, 5.594419, 5.387138, 
    5.139074, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  5.62, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  5.62, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  5.62, 5.608697, 5.600054, 5.594069, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _,
  4.38, 4.65, 4.6, 4.95, 5, 4.62, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _,
  4.38, 4.65, 4.6, 4.95, 5, 4.62, 5.594419, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _,
  4.38, 4.65, 4.6, 4.95, 5, 4.62, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _,
  4.38, 4.65, 4.6, 4.95, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _,
  4.38, 4.65, 4.6, 4.95, 5, 4.62, 5.594419, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _,
  7.72, 7.716667, 7.669908, 7.57, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _,
  7.72, 7.716667, 7.669908, 7.57, 5, 4.62, 5.594419, 5.387138, 5.139074, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  5.59, 5.531478, 5.481746, 5.440804, 5.385294, 5.3999, 5.414815, 5.397182, 
    5.340667, 5.180305, 5.233016, _, _, _, _, _, _, _, 1.96344, 1.757018, _, 
    _, _, _, _, _,
  6.08, 5.934667, 5.82, 5.736566, 5.66, 4.94, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _,
  6.08, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  6.08, 5.934667, 5.82, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _,
  6.08, 5.934667, 5.82, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _,
  6.08, 5.934667, 5.82, 5.736566, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _,
  6.08, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  6.08, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  5.6, 5.47, 5.45, 5.05, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _,
  5.6, 5.47, 5.45, 5.05, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _,
  5.6, 5.47, 5.45, 5.05, 5.66, 4.94, 5.414815, 5.397182, 5.340667, 5.180305, 
    5.233016, _, _, _, _, _, _, _, 1.96344, 1.757018, _, _, _, _, _, _,
  4.32, 4.55, 4.59, 4.66, 4.62, 4.22, 3.65, _, _, _, _, 3.93, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _,
  4.32, 4.55, 4.59, 4.66, 4.62, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _,
  5.55, 5.525886, 5.505829, 5.489829, 5.47, 5.475392, 5.482927, 5.213427, 
    4.797539, _, 3.13936, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  5.55, 5.525886, 5.505829, 5.489829, 5.47, 5.475392, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _,
  6.02, 5.963334, 5.9, 5.829134, 5.67, 5.458792, 5.2, _, 3.962494, 2.71, 
    2.06875, 1.83, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  6.02, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  6.02, 5.963334, 5.9, 5.829134, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _,
  6.02, 5.963334, 5.9, 5.829134, 5.67, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _,
  4.24, 4.37, 4.67, 4.731429, 4.59, 4.08, 3.76, 3.805, 3.85, 4.92, 5.05, 
    4.13, 4.68, 4.51, _, _, _, _, _, _, _, _, _, _, _, _,
  4.24, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  4.24, 4.37, 4.67, 4.731429, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _,
  5.49, 5.440552, 5.401989, 5.374308, 5.369231, 5.387468, 5.431084, 5.473018, 
    5.514453, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  5.49, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  5.49, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  5.49, 5.440552, 5.401989, 5.374308, 5.369231, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _,
  5.49, 5.440552, 5.401989, 5.374308, 5.369231, 5.387468, 5.431084, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  5.49, 5.440552, 5.401989, 5.374308, 5.369231, 5.387468, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  6.13, 6.252222, 6.331959, 6.205755, 6.175712, 6.15401, 6.126458, 6.097378, 
    6.01563, 5.638904, _, _, _, _, 5.038765, _, _, _, _, _, _, _, _, _, _, _,
  5.74, 5.908052, 5.958657, 5.877481, 5.444124, 4.543561, _, _, _, _, _, _, 
    _, _, _, _, _, 0.5082346, 0.5989192, 0.6816325, _, _, _, _, _, _,
  5.74, 5.908052, 5.958657, 5.877481, 5.444124, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _,
  5.74, 5.908052, 5.958657, 5.877481, 5.444124, 4.543561, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  5.74, 5.908052, 5.958657, 5.877481, 5.444124, 4.543561, _, _, _, _, _, _, 
    _, _, _, _, _, 0.5082346, 0.5989192, 0.6816325, _, _, _, _, _, _,
  5.74, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  5.74, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  4.72, 4.75, 4.76, 4.76, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _,
  4.72, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  4.72, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  4.72, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  4.72, 4.75, 4.76, 4.76, 5.444124, 4.543561, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _,
  4.72, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  4.72, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  4.72, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  4.72, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _ ;

 Oxygen_sigfigs =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  6, 6, 6, 6, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, 3, 3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, 3, 3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, 3, 3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, 3, 3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, 3, 3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, 3, 3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, 3, 3, 3, 3, 3, _, _, _, _, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, 3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, 3, 3, 3, 3, 3, _, _, _, _, 3, _, _, _, _, _, _, 2, 2, 2, _, _, _, _, _, _,
  1, 3, 3, 3, 3, 3, 3, _, 3, 3, _, _, _, 2, _, _, 2, 2, 2, 2, 2, _, _, _, _, _,
  1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, 3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, 3, 3, 3, 3, 3, 3, 3, 3, _, _, _, 3, _, _, 3, 3, 3, _, _, _, _, 3, _, 3,
  3, 3, 3, 3, 3, 3, 3, 3, 3, 3, _, _, _, 3, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, 3, 3, 3, 3, 3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, 3, 3, 3, 3, 3, 3, 3, 3, 3, _, _, _, 3, _, _, _, _, 3, 3, _, _, _, _, _, _,
  3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _,
  3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, _, _, _, 3, 3, _, _, _, _, _, _,
  3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, 3, 3, 3, 3, 3, 3, 3, 3, _, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, _, 3,
  3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, 3, 3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, 3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, 3, 3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, 3, 3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, 3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, 3, 3, 3, 3, 3, _, 3, _, 3, _, _, 3, _, _, _, 3, 3, _, _, _, _, _, _, _,
  3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _,
  1, 3, 3, 3, 3, 3, 3, _, 3, 3, _, _, _, 2, _, _, 2, 2, 2, 2, 2, _, _, _, _, _,
  1, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, 3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, 3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, 3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, 3, 3, 3, 3, 3, 3, _, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, 3, 3, 3, 3, 3, 3, _, 3, 3, _, _, _, 2, _, _, 2, 2, 2, 2, 2, _, _, _, _, _,
  1, 3, 3, 3, 3, 3, 3, _, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, 3, 3, 3, 3, 3, 3, 3, 3, 3, _, _, _, _, _, _, _, _, 3, _, _, _, _, _, _, _,
  1, 3, 3, 3, 3, 3, 3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, _, _, _, _, _, _, _, _, _, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, 3, 3, 3, 3, 3, 3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, 3, 3, 3, 3, 3, 3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, 3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, 3, 3, 3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, 3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, 3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, 3, 3, 3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, 3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, _, 3,
  1, 3, 3, 3, 3, 3, 3, _, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, 3, 3, 3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, 3, 3, 3, 3, 3, 3, _, 3, 3, 3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _,
  1, 3, 3, 3, 3, 3, 3, _, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, 3, 3, 3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, 3, 3, 3, 3, 3, 3, 3, 3, 3, _, _, _, _, _, _, _, 3, _, _, _, _, _, _, _, _,
  1, 3, 3, 3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, 3, 3, 3, 3, 3, 3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, 3, _, _, _, _, _, 3, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, 3, _, _, _, _, _, 3, _, _, _, _, _, _, _, _,
  1, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, 3, 3, 3, 3, 3, 3, 3, 3, _, 3, 3, 3, _, _, 3, 3, 3, _, _, _, _, _, _, 3,
  3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, 3, 3, 3, 3, 3, 3, 3, 3, _, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, 3, 3, 3, 3, 3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, 3, 3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, 3, 3, 3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, 3, 3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, 3, 3, 3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, 3, 3, 3, 3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, _, _, _, _, _, _, _, 3, 3, _, _, _, _, _, _,
  1, 3, 3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, _, _, _, _, _, _, _, 3, 3, _, _, _, _, _, _,
  3, 3, 3, 3, 3, 3, 3, _, _, _, _, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, 3, 3, 3, 3, 3, 3, 3, 3, _, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, 3, 3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, 3, 3, 3, 3, 3, 3, _, 3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, 3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _,
  1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, 3, 3, 3, 3, 3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, 3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, 3, 3, 3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, 3, 3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4, 4, 4, 4, 4, 4, 4, 4, 4, 4, _, _, _, _, 4, _, _, _, _, _, _, _, _, _, _, _,
  1, 3, 3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, 2, 2, 2, _, _, _, _, _, _,
  1, 3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, 3, 3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, 3, 3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, 2, 2, 2, _, _, _, _, _, _,
  1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, 3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 Oxygen_WODflag =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, _, _, _, _, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, _, _, _, _, 0, _, _, _, _, _, _, 0, 0, 0, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, 0, 0, _, _, _, 0, _, _, 0, 0, 0, 0, 0, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, 0, _, _, 0, 0, 0, _, _, _, _, 0, _, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, 0, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, 0, _, _, _, _, 0, 0, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, 0, 0, _, _, _, _, _, _,
  0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, _, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, 0,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, 0, _, 0, _, _, 0, _, _, _, 0, 0, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, 0, 0, _, _, _, 0, _, _, 0, 0, 0, 0, 0, _, _, _, _, _,
  0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, 0, 0, _, _, _, 0, _, _, 0, 0, 0, 0, 0, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, 0, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, _, _, _, _, _, _, _, _, _, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, 0,
  0, 0, 0, 0, 0, 0, 0, _, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, 6, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, 0, _, _, _, _, _, 0, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, 0, _, _, _, _, _, 0, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 9, 0, 0, 0, 0, 0, 0, 0, 0, _, 0, 0, 0, _, _, 0, 0, 0, _, _, _, _, _, _, 0,
  0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4, 4, 4, 0, 4, 4, 0, 0, 0, _, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, 0, 0, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, 0, 0, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, _, _, _, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, _, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, 0, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, 0, 0, 0, _, _, _, _, _, _,
  0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, 0, 0, 0, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 Oxygen_WODprofileflag = _, _, _, _, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 0, 
    4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0 ;

 Oxygen_Original_units =
  "ug-at/l            mmol/m3  umol/l  uM  umol/dm3",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "" ;

 Phosphate =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 0.557, 0.476, 0.542, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _,
  0.5165673, 0.4519964, 0.4519964, 0.4519964, 0.4519964, 0.4519964, 
    0.4519964, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0.5165673, 0.4519964, 0.4519964, 0.4519964, 0.4519964, 0.4519964, 
    0.4519964, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0.5165673, 0.4519964, 0.4519964, 0.4519964, 0.4519964, 0.4519964, 
    0.4519964, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0.5165673, 0.4519964, 0.4519964, 0.4519964, 0.4519964, 0.4519964, 
    0.4519964, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0.5165673, 0.4519964, 0.4519964, 0.4519964, 0.4519964, 0.4519964, 
    0.4519964, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0.5165673, 0.4519964, 0.4519964, 0.4519964, 0.4519964, 0.4519964, 
    0.4519964, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1.31138, 1.333739, 1.34691, 1.34691, 1.359309, 1.49954, _, _, _, _, 
    1.961835, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1.31138, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _,
  0.31, 0.39, 0.33, 0.41, 0.46, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _,
  0.31, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  0.31, 0.39, 0.33, 0.41, 0.46, 1.49954, _, _, _, _, 1.961835, _, _, _, _, _, 
    _, 2.801082, 3.101802, 3.385359, 1.24, 1.276744, 1.330265, 1.379, _, _,
  0.20349, 0.3182626, 0.4199, 0.5062017, 0.646, 0.7911003, 0.9044, _, 
    1.108967, 1.2597, _, _, _, 1.7765, _, _, 2.3256, 2.616299, 2.907, 3.1977, 
    3.4884, _, _, _, _, _,
  0.20349, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _,
  0.20349, 0.3182626, 0.4199, 0.5062017, 0.646, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _,
  0.20349, 0.3182626, 0.4199, 0.5062017, 0.646, 0.7911003, 0.9044, _, 
    1.108967, 1.2597, _, _, _, 1.7765, _, _, 2.3256, 2.616299, 2.907, 3.1977, 
    3.4884, 1.276744, 1.330265, 1.379, _, 1.310066,
  0.20349, 0.3182626, 0.4199, 0.5062017, 0.646, 0.7911003, 0.9044, _, 
    1.108967, 1.2597, _, _, _, 1.7765, _, _, _, _, _, _, _, _, _, _, _, _,
  0.20349, 0.3182626, 0.4199, 0.5062017, 0.646, 0.7911003, 0.9044, _, 
    1.108967, 1.2597, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0.20349, 0.3182626, 0.4199, 0.5062017, 0.646, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _,
  0.20349, 0.3182626, 0.4199, 0.5062017, 0.646, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _,
  0.20349, 0.3182626, 0.4199, 0.5062017, 0.646, 0.7911003, 0.9044, _, 
    1.108967, 1.2597, _, _, _, 1.7765, _, _, 2.3256, 2.616299, 2.907, 3.1977, 
    3.4884, 1.276744, 1.330265, 1.379, _, _,
  0.20349, 0.3182626, 0.4199, 0.5062017, 0.646, 0.7911003, 0.9044, _, 
    1.108967, 1.2597, _, _, _, 1.7765, _, _, _, _, _, _, _, _, _, _, _, _,
  0.20349, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _,
  0.25, 0.4, 0.36, 0.37, 0.37, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _,
  0.25, 0.4, 0.36, 0.37, 0.37, 0.7911003, 0.9044, _, 1.108967, 1.2597, _, _, 
    _, 1.7765, _, _, 2.3256, 2.616299, 2.907, 3.1977, 3.4884, 1.276744, 
    1.330265, 1.379, _, _,
  0.3, 0.3, 0.28, 0.41, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _,
  0.3, 0.3, 0.28, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _,
  0.3, 0.3, 0.28, 0.41, 0.37, 0.7911003, 0.9044, _, 1.108967, 1.2597, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0.3, 0.3, 0.28, 0.41, 0.37, 0.7911003, 0.9044, _, 1.108967, 1.2597, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0.3, 0.3, 0.28, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _,
  0.53, 0.53, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _,
  0.53, 0.53, 0.28, 0.41, 0.37, 0.7911003, 0.9044, _, 1.108967, 1.2597, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0.2907, 0.2956566, 0.3048322, 0.3182268, 0.3576378, 0.4120907, 0.5470413, 
    0.9846376, 1.312872, _, 1.615, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1.14, 1.14, 1.14, 1.14, 1.149, 1.149, 1.188, 1.188, 1.188, 1.227, 1.35, 
    1.269, 1.35, 1.408, 1.45, 1.417, 1.479, 1.558893, 1.65, 1.51969, 1.417, 
    1.445823, 1.473695, 1.498, _, 1.47923,
  1.14, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  1.14, 1.14, 1.14, 1.14, 1.149, 1.149, 1.188, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _,
  1.14, 1.14, 1.14, 1.14, 1.149, 1.149, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _,
  0.14, 0.19, 0.41, 0.66, 0.65, 0.639107, 0.63, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _,
  0.14, 0.19, 0.41, 0.66, 0.65, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _,
  0.14, 0.19, 0.41, 0.66, 0.65, 0.639107, 0.63, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _,
  0.14, 0.19, 0.41, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _,
  0.14, 0.19, 0.41, 0.66, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _,
  0.05, 0.19, 0.34, 0.65, 0.61, 0.63, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _,
  0.05, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  0.05, 0.19, 0.34, 0.65, 0.61, 0.63, 0.63, 1.188, 1.188, 1.227, 1.35, 1.269, 
    1.35, 1.408, 1.45, 1.417, 1.479, 1.558893, 1.65, 1.51969, 1.417, 
    1.445823, 1.473695, 1.498, _, _,
  0.05, 0.19, 0.34, 0.65, 0.61, 0.63, 0.63, 1.188, 1.188, 1.227, 1.35, 1.269, 
    1.35, 1.408, 1.45, _, _, _, _, _, _, _, _, _, _, _,
  0.05, 0.19, 0.34, 0.65, 0.61, 0.63, 0.63, 1.188, 1.188, 1.227, 1.35, 1.269, 
    1.35, 1.408, 1.45, 1.417, 1.479, 1.558893, 1.65, 1.51969, 1.417, _, _, _, 
    _, _,
  0.53, 0.63, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _,
  0.53, 0.63, 0.34, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _,
  0.53, 0.63, 0.34, 0.65, 0.61, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _,
  0.53, 0.63, 0.34, 0.65, 0.61, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _,
  0.53, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  0.53, 0.63, 0.34, 0.65, 0.61, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _,
  0.53, 0.63, 0.34, 0.65, 0.61, 0.63, 0.63, 1.188, 1.188, 1.227, 1.35, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _,
  0.53, 0.63, 0.34, 0.65, 0.61, 0.63, 0.63, 1.188, 1.188, 1.227, 1.35, 1.269, 
    1.35, 1.408, 1.45, 1.417, 1.479, 1.558893, 1.65, 1.51969, 1.417, 
    1.445823, 1.473695, 1.498, _, _,
  0.1, 0.6, 0.71, 0.68, 0.63, 0.6676785, 0.7, 0.714192, 0.73, 0.77, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _,
  0.1, 0.6, 0.71, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _,
  0.6, 0.63, 0.61, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _,
  0.62, 0.55, 0.55, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _,
  0.62, 0.55, 0.55, 0.68, 0.63, 0.6676785, 0.7, 0.714192, 0.73, 0.77, 1.35, 
    1.269, 1.35, 1.408, 1.45, 1.417, 1.479, 1.558893, 1.65, 1.51969, 1.417, 
    1.445823, 1.473695, 1.498, _, _,
  0.62, 0.55, 0.55, 0.68, 0.63, 0.6676785, 0.7, 0.714192, 0.73, 0.77, 1.35, 
    1.269, 1.35, 1.408, 1.45, 1.417, _, _, _, _, _, _, _, _, _, _,
  0.09, 0.58, 0.66, 0.61, 0.68, 0.65652, 0.65, 0.7058163, 0.75, 0.8, _, 0.8, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0.09, 0.58, 0.66, 0.61, 0.68, 0.65652, 0.65, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _,
  0.09, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  0.09, 0.58, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _,
  0.09, 0.58, 0.66, 0.61, 0.68, 0.65652, 0.65, 0.7058163, 0.75, 0.8, _, 0.8, 
    1.35, 1.408, 1.45, 1.417, _, _, _, _, _, _, _, _, _, _,
  0.6, 0.55, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _,
  0.6, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  0.07, 0.05, 0.54, 0.51, 0.56, 0.6294, 0.7, 0.7656757, 0.82, 0.82, _, 0.784, 
    0.7, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0.6, 0.61, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _,
  0.6, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  0.27455, 0.2670104, 0.2562029, 0.2421274, 0.2030548, 0.1370363, 0.2614298, 
    0.488659, 0.7309672, 1.097384, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  0.27455, 0.2670104, 0.2562029, 0.2421274, 0.2030548, 0.1370363, 0.2614298, 
    0.488659, 0.7309672, 1.097384, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  0.27455, 0.2670104, 0.2562029, 0.2421274, 0.2030548, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0.27455, 0.2670104, 0.2562029, 0.2421274, 0.2030548, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0.17, 0.15, 0.2636364, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _,
  0.37, 0.26, 0.35, 0.32, 0.35, 0.32, 1.39, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _,
  0.37, 0.26, 0.35, 0.32, 0.35, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _,
  0.37, 0.26, 0.35, 0.32, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _,
  0.49, 0.61, 0.5766667, 0.5433334, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _,
  0.49, 0.61, 0.5766667, 0.5433334, _, 0.32, 1.39, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _,
  0.02, 0.06, 0.59, 0.59, 0.58, 0.5965704, 0.64, 0.69625, 0.77, _, _, _, 
    0.78, 0.6875556, 0.54, _, _, _, _, _, _, _, _, _, _, _,
  0.02, 0.06, 0.59, 0.59, 0.58, 0.5965704, 0.64, 0.69625, 0.77, _, _, _, 
    0.78, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1.107, 1.078, 1.078, 1.078, 1.078, 1.03, 1.14, 1.079098, 1.049, 1.117, 
    1.178, 1.217, 1.198, 1.198, 1.198, 1.259, 1.198, 1.198, 1.198, 1.21384, 
    1.24, 1.276744, 1.330265, 1.379, _, 1.310066,
  0.25194, 0.3570227, 0.4522, 0.5360556, 0.6783, 0.8234002, 0.9367, _, 
    1.141267, 1.292, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0.25194, 0.3570227, 0.4522, 0.5360556, 0.6783, 0.8234002, 0.9367, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0.25194, 0.3570227, 0.4522, 0.5360556, 0.6783, 0.8234002, 0.9367, _, 
    1.141267, 1.292, 1.178, 1.217, 1.198, 1.198, _, _, _, _, _, _, _, _, _, 
    _, _, _,
  0.25194, 0.3570227, 0.4522, 0.5360556, 0.6783, 0.8234002, 0.9367, _, 
    1.141267, 1.292, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0.4, 0.53, 0.44, 0.44, 0.43, 0.43, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _,
  0.4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  0.4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  0.4, 0.53, 0.44, 0.44, 0.43, 0.43, _, _, 1.141267, 1.292, 1.178, 1.217, 
    1.198, 1.198, 1.198, 1.259, 1.198, 1.198, 1.198, 1.21384, 1.24, 1.276744, 
    1.330265, 1.379, _, _,
  0.4, 0.53, 0.44, 0.44, 0.43, 0.43, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _,
  0.4, 0.53, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _,
  0.4, 0.53, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _,
  0.4, 0.53, 0.44, 0.44, 0.43, 0.43, _, _, 1.141267, 1.292, 1.178, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _,
  0.08, 0.19, 0.56, 0.54, 0.56, 0.6097453, 0.67, 0.67, 0.67, 0.64, _, 
    0.6701316, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0.08, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  0.08, 0.19, 0.56, 0.54, 0.56, 0.6097453, 0.67, 0.67, 0.67, 0.64, _, 
    0.6701316, 1.198, 1.198, 1.198, 1.259, 1.198, 1.198, 1.198, 1.21384, 
    1.24, 1.276744, 1.330265, 1.379, _, _,
  0.08, 0.19, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _,
  0.08, 0.19, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _,
  0.08, 0.19, 0.56, 0.54, 0.56, 0.6097453, 0.67, 0.67, 0.67, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _,
  0.08, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  0.08, 0.19, 0.56, 0.54, 0.56, 0.6097453, 0.67, 0.67, 0.67, 0.64, _, 
    0.6701316, 1.198, 1.198, 1.198, 1.259, 1.198, 1.198, 1.198, 1.21384, 
    1.24, 1.276744, 1.330265, 1.379, _, _,
  0.15, 0.1418182, 0.1743899, 0.24, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _,
  0.15, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  0.15, 0.1418182, 0.1743899, 0.24, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _,
  0.15, 0.1418182, 0.1743899, 0.24, 0.56, 0.6097453, 0.67, 0.67, 0.67, 0.64, 
    _, 0.6701316, 1.198, 1.198, 1.198, 1.259, 1.198, 1.198, 1.198, 1.21384, 
    1.24, 1.276744, 1.330265, 1.379, _, 1.310066,
  0.15, 0.1418182, 0.1743899, 0.24, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _,
  0.31008, 0.2751771, 0.2512066, 0.2676862, 0.2452916, 0.3178998, 0.4456995, 
    0.5978347, 0.8105975, _, 1.648351, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  0.18, 0.24, 0.53, 0.53, 0.51, 0.5254405, 0.54, 0.5528921, 0.56, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _,
  0.18, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  0.18, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  0.18, 0.24, 0.53, 0.53, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _,
  0.15, 0.1418182, 0.1609646, 0.223959, 0.3159886, 0.42, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _,
  0.15, 0.1418182, 0.1609646, 0.223959, 0.3159886, 0.42, 0.54, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0.26, 0.4, 0.4, 0.54, 0.53, 0.53, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _,
  0.26, 0.4, 0.4, 0.54, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _,
  0.26, 0.4, 0.4, 0.54, 0.53, 0.53, 0.54, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _,
  0.26, 0.4, 0.4, 0.54, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _,
  0.26, 0.4, 0.4, 0.54, 0.53, 0.53, 0.54, 0.5528921, 0.56, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _,
  0.26, 0.4, 0.4, 0.54, 0.53, 0.53, 0.54, 0.5528921, 0.56, _, 1.648351, _, _, 
    _, _, _, _, _, _, _, 1.24, 1.276744, 1.330265, 1.379, _, _,
  0.3553, 0.4608133, 0.5491, 0.5993958, 0.7106, 0.8721, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _,
  0.3553, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _,
  0.3553, 0.4608133, 0.5491, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _,
  0.3553, 0.4608133, 0.5491, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _,
  0.18, 0.26, 0.38, 0.46, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _,
  0.18, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  0.18, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  0.18, 0.26, 0.38, 0.46, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _,
  0.18, 0.26, 0.38, 0.46, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _,
  0.18, 0.26, 0.38, 0.46, 0.7106, 0.8721, 0.54, 0.5528921, 0.56, _, 1.648351, 
    _, _, _, _, _, _, _, _, _, 1.24, 1.276744, 1.330265, 1.379, _, _,
  0.15, 0.1572, 0.1730118, 0.2015636, 0.3373979, 0.462964, _, 0.8528858, _, 
    1.02, 1.072391, 1.112246, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0.67, 0.7, 0.62, 0.59, 0.45, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _,
  0.4522, 0.428733, 0.4105396, 0.3976196, 0.3876, 0.4205592, 0.4603345, 
    0.7624305, 1.056452, _, 1.913817, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  0.4522, 0.428733, 0.4105396, 0.3976196, 0.3876, 0.4205592, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0.4522, 0.428733, 0.4105396, 0.3976196, 0.3876, 0.4205592, 0.4603345, 
    0.7624305, 1.056452, _, 1.913817, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  0.4522, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _,
  0.4522, 0.428733, 0.4105396, 0.3976196, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _,
  0.4522, 0.428733, 0.4105396, 0.3976196, 0.3876, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _,
  0.14, 0.14, 0.1507069, 0.1766394, 0.27, 0.46, 0.63, 0.615, 0.6, 1.133447, 
    1.15913, 1.19135, 1.423645, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0.14, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  0.14, 0.14, 0.1507069, 0.1766394, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _,
  0.14, 0.14, 0.1507069, 0.1766394, 0.27, 0.46, 0.63, 0.615, 0.6, 1.133447, 
    1.15913, 1.19135, 1.423645, _, _, _, _, _, _, _, 1.24, 1.276744, _, _, _, _,
  0.14, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  0.14, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  0.14, 0.14, 0.1507069, 0.1766394, 0.27, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _,
  0.14, 0.14, 0.1507069, 0.1766394, 0.27, 0.46, 0.63, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _,
  0.14, 0.14, 0.1507069, 0.1766394, 0.27, 0.46, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _,
  0.14, 0.14, 0.1507069, 0.1766394, 0.27, 0.46, 0.63, 0.615, 0.6, 1.133447, 
    1.15913, 1.19135, 1.423645, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0.23256, 0.397553, 0.5283017, 0.6072736, 0.7293423, 0.8731752, _, _, _, _, 
    _, _, _, _, _, _, _, 2.801082, 3.101802, 3.385359, _, _, _, _, _, _,
  0.23256, 0.397553, 0.5283017, 0.6072736, 0.7293423, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _,
  0.23256, 0.397553, 0.5283017, 0.6072736, 0.7293423, 0.8731752, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0.23256, 0.397553, 0.5283017, 0.6072736, 0.7293423, 0.8731752, _, _, _, _, 
    _, _, _, _, _, _, _, 2.801082, 3.101802, 3.385359, 1.24, 1.276744, 
    1.330265, 1.379, _, _,
  0.55, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  0.66, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  0.66, 0.397553, 0.5283017, 0.6072736, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _,
  0.67, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  0.67, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  0.51, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  0.51, 0.397553, 0.5283017, 0.6072736, 0.7293423, 0.8731752, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0.5, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  0.74, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  0.55, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  0.49, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _ ;

 Phosphate_sigfigs =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4, 4, 4, 4, 4, 4, 4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4, 4, 4, 4, 4, 4, 4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4, 4, 4, 4, 4, 4, 4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4, 4, 4, 4, 4, 4, 4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4, 4, 4, 4, 4, 4, 4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4, 4, 4, 4, 4, 4, 4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, 3, 3, 3, 3, 3, _, _, _, _, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, 2, 3, _, _, _, _, 3, _, _, _, _, _, _, 3, 3, 3, 4, 4, 4, 4, _, _,
  1, 2, 3, 3, 3, 3, 3, _, 3, 3, _, _, _, 3, _, _, 3, 3, 3, 3, 4, _, _, _, _, _,
  1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, 2, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, 2, 3, 3, 3, 3, 3, _, 3, 3, _, _, _, 3, _, _, 3, 3, 3, 3, 4, 4, 4, 4, _, 4,
  1, 2, 3, 3, 3, 3, 3, _, 3, 3, _, _, _, 3, _, _, _, _, _, _, _, _, _, _, _, _,
  1, 2, 3, 3, 3, 3, 3, _, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, 2, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, 2, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, 2, 3, 3, 3, 3, 3, _, 3, 3, _, _, _, 3, _, _, 3, 3, 3, 3, 4, 4, 4, 4, _, _,
  1, 2, 3, 3, 3, 3, 3, _, 3, 3, _, _, _, 3, _, _, _, _, _, _, _, _, _, _, _, _,
  1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, 2, 3, 3, _, 3, 3, _, _, _, 3, _, _, 3, 3, 3, 3, 4, 4, 4, 4, _, _,
  2, 2, 2, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, 2, 3, 3, _, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, 2, 3, 3, _, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, 2, 3, 3, _, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, 2, 2, 2, 3, 3, 2, 2, 3, _, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, _, 4,
  4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4, 4, 4, 4, 4, 4, 4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4, 4, 4, 4, 4, 4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, 2, 2, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, 2, 2, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, 2, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, 2, 2, 2, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, _, _,
  2, 2, 2, 2, 2, 2, 2, 4, 4, 4, 4, 4, 4, 4, 4, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, 2, 2, 2, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, _, _, _, _, _,
  2, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, 2, 2, 2, 4, 4, 4, 4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, 2, 2, 2, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, _, _,
  2, 2, 2, 2, 2, 2, 2, 2, 2, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, _, _,
  2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 4, 4, 4, 4, 4, 4, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, 2, 2, 2, 2, 2, 2, _, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, 2, 2, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, 2, 2, 2, 2, 2, 2, _, 2, 4, 4, 4, 4, _, _, _, _, _, _, _, _, _, _,
  2, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, 2, 2, 2, 2, 2, 2, _, 2, 2, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, 2, 2, 2, 2, 2, 2, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, 2, 2, 2, 2, 2, 2, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, 2, 2, 2, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, 2, 2, 2, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, 2, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, 2, 2, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, _, 2, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, 2, 2, 2, 2, 2, _, _, _, 2, 2, 2, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, 2, 2, 2, 2, 2, _, _, _, 2, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, _, 4,
  1, 2, 3, 3, 3, 3, 3, _, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, 2, 3, 3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, 2, 3, 3, 3, 3, 3, _, 3, 3, 4, 4, 4, 4, _, _, _, _, _, _, _, _, _, _, _, _,
  1, 2, 3, 3, 3, 3, 3, _, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, 2, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, 2, 2, _, _, 3, 3, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, _, _,
  2, 2, 2, 2, 2, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, 2, 2, _, _, 3, 3, 4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, 2, 2, 2, 2, 2, 2, _, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, 2, 2, 2, 2, 2, 2, _, 2, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, _, _,
  2, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, 2, 2, 2, 2, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, 2, 2, 2, 2, 2, 2, _, 2, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, _, _,
  1, 2, 2, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, 2, 2, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, 2, 2, 2, 2, 2, 2, 2, 2, 2, _, 2, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, _, 4,
  1, 2, 2, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, 2, 2, 2, 2, 2, 3, 3, 2, _, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, 2, 2, 2, 2, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, 2, 2, 2, 2, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, 2, 2, 2, 2, 2, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, 2, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, 2, 2, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, 2, 2, 2, 2, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, 2, 2, 2, 2, 2, _, 3, _, _, _, _, _, _, _, _, _, 4, 4, 4, 4, _, _,
  1, 3, 3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, 3, 3, 2, 2, 2, _, 3, _, _, _, _, _, _, _, _, _, 4, 4, 4, 4, _, _,
  1, 2, 2, 2, 2, 2, _, 2, _, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, 3, 3, 3, 3, 3, 2, 2, 3, _, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, 3, 3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, 3, 3, 3, 3, 3, 2, 2, 3, _, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, 3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, 2, 2, 2, 2, 2, 2, 2, 2, 3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, 2, 2, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, 2, 2, 2, 2, 2, 2, 2, 2, 3, 3, 3, 3, _, _, _, _, _, _, _, 4, 4, _, _, _, _,
  1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, 2, 2, 2, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, 2, 2, 2, 2, 2, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, 2, 2, 2, 2, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, 2, 2, 2, 2, 2, 2, 2, 2, 3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, 2, 3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, 3, 3, 3, _, _, _, _, _, _,
  1, 2, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, 2, 3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, 2, 3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, 3, 3, 3, 4, 4, 4, 4, _, _,
  1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, 2, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, 2, 3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 Phosphate_WODflag =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, _, _, _, _, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, _, _, _, _, 0, _, _, _, _, _, _, 0, 0, 0, 0, 0, 0, 0, _, _,
  0, 0, 0, 0, 0, 0, 0, _, 0, 6, _, _, _, 6, _, _, 6, 1, 1, 0, 0, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, 0, 0, _, _, _, 0, _, _, 0, 0, 0, 0, 0, 0, 0, 0, _, 0,
  0, 0, 0, 0, 0, 0, 0, _, 0, 0, _, _, _, 0, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, 0, 0, _, _, _, 0, _, _, 0, 0, 0, 0, 0, 0, 0, 0, _, _,
  0, 0, 0, 0, 0, 0, 0, _, 0, 0, _, _, _, 0, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, 0, 0, _, _, _, 0, _, _, 0, 0, 0, 0, 0, 0, 0, 0, _, _,
  0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, _, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 3, 3, 0, 0, 3, 3, _, 7,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _,
  0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _,
  0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, _, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, 0, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, 0,
  0, 0, 0, 0, 0, 0, 0, _, 0, 6, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, _, _, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _,
  0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, _, _, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _,
  0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _,
  0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, 0,
  0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, _, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, _, 0, _, _, _, _, _, _, _, _, _, 0, 0, 0, 0, _, _,
  0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, _, 0, _, _, _, _, _, _, _, _, _, 0, 0, 0, 0, _, _,
  0, 0, 0, 0, 0, 0, _, 0, _, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, _, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, _, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, 0, 0, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, 0, 0, 0, _, _, _, _, _, _,
  0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, 0, 0, 0, 0, 0, 0, 0, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 Phosphate_WODprofileflag = _, _, _, _, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 Phosphate_Original_units =
  "\"ug/l\"    Alternate Nutrient Conversion (use instead of #36)",
  "\"ug/l\"    Alternate Nutrient Conversion (use instead of #36)",
  "ug/l               mg/m3    ppb     g/1000m3",
  "\"ug/l\"    Alternate Nutrient Conversion (use instead of #36)",
  "\"ug/l\"    Alternate Nutrient Conversion (use instead of #36)",
  "ug/l               mg/m3    ppb     g/1000m3",
  "\"ug/l\"    Alternate Nutrient Conversion (use instead of #36)",
  "ug/l               mg/m3    ppb     g/1000m3",
  "\"ug/l\"    Alternate Nutrient Conversion (use instead of #36)",
  "ug/l               mg/m3    ppb     g/1000m3",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "" ;

 TotalPhos =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0.07, 0.0478836, 0.03, 0.02136364, 0.03169274, 0.11, 0.283451, _, 
    0.4395986, _, 0.3840765, _, _, 0.6772242, _, _, _, 0.7215907, 0.656701, 
    _, _, _, _, _, _, _,
  0.07, 0.0478836, 0.03, 0.02136364, 0.03169274, 0.11, 0.283451, _, 
    0.4395986, _, 0.3840765, _, _, 0.6772242, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  0.07, 0.0478836, 0.03, 0.02136364, 0.03169274, 0.11, 0.283451, _, 
    0.4395986, _, 0.3840765, _, _, 0.6772242, _, _, _, 0.7215907, 0.656701, 
    _, _, _, _, _, _, _,
  0.07, 0.0478836, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _,
  0.07, 0.0478836, 0.03, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _,
  0.07, 0.0478836, 0.03, 0.02136364, 0.03169274, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _,
  0.07, 0.0478836, 0.03, 0.02136364, 0.03169274, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _,
  0.07, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  0.07, 0.0478836, 0.03, 0.02136364, 0.03169274, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _,
  0.07, 0.0478836, 0.03, 0.02136364, 0.03169274, 0.11, 0.283451, _, 
    0.4395986, _, 0.3840765, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0.07, 0.0478836, 0.03, 0.02136364, 0.03169274, 0.11, 0.283451, _, 
    0.4395986, _, 0.3840765, _, _, 0.6772242, _, _, _, 0.7215907, 0.656701, 
    _, _, _, _, _, _, _,
  0.07, 0.0478836, 0.03, 0.02136364, 0.03169274, 0.11, 0.283451, _, 
    0.4395986, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0.07, 0.0478836, 0.03, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _,
  0.07, 0.0478836, 0.03, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _,
  0.07, 0.0478836, 0.03, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _,
  0.07, 0.0478836, 0.03, 0.02136364, 0.03169274, 0.11, 0.283451, _, 
    0.4395986, _, 0.3840765, _, _, 0.6772242, _, _, _, 0.7215907, 0.656701, 
    _, _, _, _, _, _, _,
  0.07, 0.0478836, 0.03, 0.02136364, 0.03169274, 0.11, 0.283451, _, 
    0.4395986, _, 0.3840765, _, _, 0.6772242, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  0.07, 0.0478836, 0.03, 0.02136364, 0.03169274, 0.11, 0.283451, _, 
    0.4395986, _, 0.3840765, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0.07, 0.0478836, 0.03, 0.02136364, 0.03169274, 0.11, 0.283451, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0.07, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  0.07, 0.0478836, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _,
  0.07, 0.0478836, 0.03, 0.02136364, 0.03169274, 0.11, 0.283451, _, 
    0.4395986, _, 0.3840765, _, _, 0.6772242, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  0.07, 0.0478836, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _,
  0.07, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  0.07, 0.0478836, 0.03, 0.02136364, 0.03169274, 0.11, 0.283451, _, 
    0.4395986, _, 0.3840765, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0.07, 0.0478836, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _,
  0.07, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  0.07, 0.0478836, 0.03, 0.02136364, 0.03169274, 0.11, 0.283451, _, 
    0.4395986, _, 0.3840765, _, _, 0.6772242, _, _, _, 0.7215907, 0.656701, 
    _, _, _, _, _, _, _,
  0.07, 0.0478836, 0.03, 0.02136364, 0.03169274, 0.11, 0.283451, _, 
    0.4395986, _, 0.3840765, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0.07, 0.0478836, 0.03, 0.02136364, 0.03169274, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _,
  0.07, 0.0478836, 0.03, 0.02136364, 0.03169274, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _,
  0.07, 0.0478836, 0.03, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _,
  0.07, 0.0478836, 0.03, 0.02136364, 0.03169274, 0.11, 0.283451, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0.07, 0.0478836, 0.03, 0.02136364, 0.03169274, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _,
  0.07, 0.0478836, 0.03, 0.02136364, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _,
  0.07, 0.0478836, 0.03, 0.02136364, 0.03169274, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _,
  0.07, 0.0478836, 0.03, 0.02136364, 0.03169274, 0.11, 0.283451, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0.07, 0.0478836, 0.03, 0.02136364, 0.03169274, 0.11, 0.283451, _, 
    0.4395986, _, 0.3840765, _, _, 0.6772242, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  0.07, 0.0478836, 0.03, 0.02136364, 0.03169274, 0.11, 0.283451, _, 
    0.4395986, _, 0.3840765, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0.07, 0.0478836, 0.03, 0.02136364, 0.03169274, 0.11, 0.283451, _, 
    0.4395986, _, 0.3840765, _, _, 0.6772242, _, _, _, 0.7215907, 0.656701, 
    _, _, _, _, _, _, _,
  0.07, 0.0478836, 0.03, 0.02136364, 0.03169274, 0.11, 0.283451, _, 
    0.4395986, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0.07, 0.0478836, 0.03, 0.02136364, 0.03169274, 0.11, 0.283451, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0.07, 0.0478836, 0.03, 0.02136364, 0.03169274, 0.11, 0.283451, _, 
    0.4395986, _, 0.3840765, _, _, 0.6772242, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  0.07, 0.0478836, 0.03, 0.02136364, 0.03169274, 0.11, 0.283451, _, 
    0.4395986, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0.07, 0.0478836, 0.03, 0.02136364, 0.03169274, 0.11, 0.283451, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0.07, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  0.07, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  0.07, 0.0478836, 0.03, 0.02136364, 0.03169274, 0.11, 0.283451, _, 
    0.4395986, _, 0.3840765, _, _, 0.6772242, _, _, _, 0.7215907, 0.656701, 
    _, _, _, _, _, _, _,
  0.07, 0.0478836, 0.03, 0.02136364, 0.03169274, 0.11, 0.283451, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0.07, 0.0478836, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _,
  0.07, 0.0478836, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _,
  0.07, 0.0478836, 0.03, 0.02136364, 0.03169274, 0.11, 0.283451, _, 
    0.4395986, _, 0.3840765, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0.07, 0.0478836, 0.03, 0.02136364, 0.03169274, 0.11, 0.283451, _, 
    0.4395986, _, 0.3840765, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0.07, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  0.07, 0.0478836, 0.03, 0.02136364, 0.03169274, 0.11, 0.283451, _, 
    0.4395986, _, 0.3840765, _, _, 0.6772242, _, _, _, 0.7215907, 0.656701, 
    _, _, _, _, _, _, _,
  0.07, 0.0478836, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _,
  0.07, 0.0478836, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _,
  0.07, 0.0478836, 0.03, 0.02136364, 0.03169274, 0.11, 0.283451, _, 
    0.4395986, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0.07, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  0.07, 0.0478836, 0.03, 0.02136364, 0.03169274, 0.11, 0.283451, _, 
    0.4395986, _, 0.3840765, _, _, 0.6772242, _, _, _, 0.7215907, 0.656701, 
    _, _, _, _, _, _, _,
  0.07, 0.0478836, 0.03, 0.02136364, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _,
  0.07, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  0.07, 0.0478836, 0.03, 0.02136364, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _,
  0.07, 0.0478836, 0.03, 0.02136364, 0.03169274, 0.11, 0.283451, _, 
    0.4395986, _, 0.3840765, _, _, 0.6772242, _, _, _, 0.7215907, 0.656701, 
    _, _, _, _, _, _, _,
  0.07, 0.0478836, 0.03, 0.02136364, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _,
  0.07, 0.0478836, 0.03, 0.02136364, 0.03169274, 0.11, 0.283451, _, 
    0.4395986, _, 0.3840765, _, _, 0.6772242, _, _, _, 0.7215907, 0.656701, 
    _, _, _, _, _, _, _,
  0.07, 0.0478836, 0.03, 0.02136364, 0.03169274, 0.11, 0.283451, _, 
    0.4395986, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0.07, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  0.07, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  0.07, 0.0478836, 0.03, 0.02136364, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _,
  0.07, 0.0478836, 0.03, 0.02136364, 0.03169274, 0.11, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _,
  0.07, 0.0478836, 0.03, 0.02136364, 0.03169274, 0.11, 0.283451, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0.07, 0.0478836, 0.03, 0.02136364, 0.03169274, 0.11, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _,
  0.07, 0.0478836, 0.03, 0.02136364, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _,
  0.07, 0.0478836, 0.03, 0.02136364, 0.03169274, 0.11, 0.283451, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0.07, 0.0478836, 0.03, 0.02136364, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _,
  0.07, 0.0478836, 0.03, 0.02136364, 0.03169274, 0.11, 0.283451, _, 
    0.4395986, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0.07, 0.0478836, 0.03, 0.02136364, 0.03169274, 0.11, 0.283451, _, 
    0.4395986, _, 0.3840765, _, _, 0.6772242, _, _, _, 0.7215907, 0.656701, 
    _, _, _, _, _, _, _,
  0.07, 0.0478836, 0.03, 0.02136364, 0.03169274, 0.11, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _,
  0.07, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  0.07, 0.0478836, 0.03, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _,
  0.07, 0.0478836, 0.03, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _,
  0.07, 0.0478836, 0.03, 0.02136364, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _,
  0.07, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  0.07, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  0.07, 0.0478836, 0.03, 0.02136364, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _,
  0.07, 0.0478836, 0.03, 0.02136364, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _,
  0.07, 0.0478836, 0.03, 0.02136364, 0.03169274, 0.11, 0.283451, _, 
    0.4395986, _, 0.3840765, _, _, 0.6772242, _, _, _, 0.7215907, 0.656701, 
    _, _, _, _, _, _, _,
  0.07, 0.0478836, 0.03, 0.02136364, 0.03169274, 0.11, 0.283451, _, 
    0.4395986, _, 0.3840765, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0.07, 0.0478836, 0.03, 0.02136364, 0.03169274, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _,
  0.07, 0.0478836, 0.03, 0.02136364, 0.03169274, 0.11, 0.283451, _, 
    0.4395986, _, 0.3840765, _, _, 0.6772242, _, _, _, 0.7215907, 0.656701, 
    _, _, _, _, _, _, _,
  0.07, 0.0478836, 0.03, 0.02136364, 0.03169274, 0.11, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _,
  0.07, 0.0478836, 0.03, 0.02136364, 0.03169274, 0.11, 0.283451, _, 
    0.4395986, _, 0.3840765, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0.07, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  0.07, 0.0478836, 0.03, 0.02136364, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _,
  0.07, 0.0478836, 0.03, 0.02136364, 0.03169274, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _,
  0.07, 0.0478836, 0.03, 0.02136364, 0.03169274, 0.11, 0.283451, _, 
    0.4395986, _, 0.3840765, _, _, 0.6772242, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  0.07, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  0.07, 0.0478836, 0.03, 0.02136364, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _,
  0.07, 0.0478836, 0.03, 0.02136364, 0.03169274, 0.11, 0.283451, _, 
    0.4395986, _, 0.3840765, _, _, 0.6772242, _, _, _, 0.7215907, 0.656701, 
    _, _, _, _, _, _, _,
  0.07, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  0.07, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  0.07, 0.0478836, 0.03, 0.02136364, 0.03169274, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _,
  0.07, 0.0478836, 0.03, 0.02136364, 0.03169274, 0.11, 0.283451, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0.07, 0.0478836, 0.03, 0.02136364, 0.03169274, 0.11, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _,
  0.07, 0.0478836, 0.03, 0.02136364, 0.03169274, 0.11, 0.283451, _, 
    0.4395986, _, 0.3840765, _, _, 0.6772242, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  0.07, 0.0478836, 0.03, 0.02136364, 0.03169274, 0.11, 0.283451, _, 
    0.4395986, _, 0.3840765, _, _, 0.6772242, _, _, _, 0.7215907, 0.656701, 
    _, _, _, _, _, _, _,
  0.07, 0.0478836, 0.03, 0.02136364, 0.03169274, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _,
  0.07, 0.0478836, 0.03, 0.02136364, 0.03169274, 0.11, 0.283451, _, 
    0.4395986, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0.07, 0.0478836, 0.03, 0.02136364, 0.03169274, 0.11, 0.283451, _, 
    0.4395986, _, 0.3840765, _, _, 0.6772242, _, _, _, 0.7215907, 0.656701, 
    _, _, _, _, _, _, _,
  0.07, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  0.07, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  0.07, 0.0478836, 0.03, 0.02136364, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _,
  0.07, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  0.07, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  0.07, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  0.07, 0.0478836, 0.03, 0.02136364, 0.03169274, 0.11, 0.283451, _, 
    0.4395986, _, 0.3840765, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0.07, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  0.07, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  0.07, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  0.07, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _ ;

 TotalPhos_sigfigs =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, 2, 2, 2, _, 2, _, 2, _, _, 2, _, _, _, 2, 2, _, _, _, _, _, _, _,
  2, 2, 2, 2, 2, 2, 2, _, 2, _, 2, _, _, 2, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, 2, 2, 2, _, 2, _, 2, _, _, 2, _, _, _, 2, 2, _, _, _, _, _, _, _,
  2, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, 2, 2, 2, _, 2, _, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, 2, 2, 2, _, 2, _, 2, _, _, 2, _, _, _, 2, 2, _, _, _, _, _, _, _,
  2, 2, 2, 2, 2, 2, 2, _, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, 2, 2, 2, _, 2, _, 2, _, _, 2, _, _, _, 2, 2, _, _, _, _, _, _, _,
  2, 2, 2, 2, 2, 2, 2, _, 2, _, 2, _, _, 2, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, 2, 2, 2, _, 2, _, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, 2, 2, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, 2, 2, 2, _, 2, _, 2, _, _, 2, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, 2, 2, 2, _, 2, _, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, 2, 2, 2, _, 2, _, 2, _, _, 2, _, _, _, 2, 2, _, _, _, _, _, _, _,
  2, 2, 2, 2, 2, 2, 2, _, 2, _, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, 2, 2, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, 2, 2, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, 2, 2, 2, _, 2, _, 2, _, _, 2, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, 2, 2, 2, _, 2, _, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, 2, 2, 2, _, 2, _, 2, _, _, 2, _, _, _, 2, 2, _, _, _, _, _, _, _,
  2, 2, 2, 2, 2, 2, 2, _, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, 2, 2, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, 2, 2, 2, _, 2, _, 2, _, _, 2, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, 2, 2, 2, _, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, 2, 2, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, 2, 2, 2, _, 2, _, 2, _, _, 2, _, _, _, 2, 2, _, _, _, _, _, _, _,
  2, 2, 2, 2, 2, 2, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, 2, 2, 2, _, 2, _, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, 2, 2, 2, _, 2, _, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, 2, 2, 2, _, 2, _, 2, _, _, 2, _, _, _, 2, 2, _, _, _, _, _, _, _,
  2, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, 2, 2, 2, _, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, 2, 2, 2, _, 2, _, 2, _, _, 2, _, _, _, 2, 2, _, _, _, _, _, _, _,
  2, 2, 2, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, 2, 2, 2, _, 2, _, 2, _, _, 2, _, _, _, 2, 2, _, _, _, _, _, _, _,
  2, 2, 2, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, 2, 2, 2, _, 2, _, 2, _, _, 2, _, _, _, 2, 2, _, _, _, _, _, _, _,
  2, 2, 2, 2, 2, 2, 2, _, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, 2, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, 2, 2, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, 2, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, 2, 2, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, 2, 2, 2, _, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, 2, 2, 2, _, 2, _, 2, _, _, 2, _, _, _, 2, 2, _, _, _, _, _, _, _,
  2, 2, 2, 2, 2, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, 2, 2, 2, _, 2, _, 2, _, _, 2, _, _, _, 2, 2, _, _, _, _, _, _, _,
  2, 2, 2, 2, 2, 2, 2, _, 2, _, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, 2, 2, 2, _, 2, _, 2, _, _, 2, _, _, _, 2, 2, _, _, _, _, _, _, _,
  2, 2, 2, 2, 2, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, 2, 2, 2, _, 2, _, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, 2, 2, 2, _, 2, _, 2, _, _, 2, _, _, _, _, _, _, _, _, _, _, _, _,
  2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, 2, 2, 2, _, 2, _, 2, _, _, 2, _, _, _, 2, 2, _, _, _, _, _, _, _,
  2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, 2, 2, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, 2, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, 2, 2, 2, _, 2, _, 2, _, _, 2, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, 2, 2, 2, _, 2, _, 2, _, _, 2, _, _, _, 2, 2, _, _, _, _, _, _, _,
  2, 2, 2, 2, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, 2, 2, 2, _, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, 2, 2, 2, _, 2, _, 2, _, _, 2, _, _, _, 2, 2, _, _, _, _, _, _, _,
  2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, 2, 2, 2, _, 2, _, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 TotalPhos_WODflag =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, 0, _, 0, _, _, 0, _, _, _, 0, 0, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, 0, _, 0, _, _, 0, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, 0, _, 0, _, _, 0, _, _, _, 0, 0, _, _, _, _, _, _, _,
  0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, 0, _, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, 0, _, 0, _, _, 0, _, _, _, 0, 0, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, 0, _, 0, _, _, 0, _, _, _, 0, 0, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, 0, _, 0, _, _, 0, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, 0, _, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, 0, _, 0, _, _, 0, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, 0, _, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, 0, _, 0, _, _, 0, _, _, _, 0, 0, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, 0, _, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, 0, _, 0, _, _, 0, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, 0, _, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, 0, _, 0, _, _, 0, _, _, _, 0, 0, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, 0, _, 0, _, _, 0, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, 0, _, 0, _, _, 0, _, _, _, 0, 0, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, 0, _, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, 0, _, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, 0, _, 0, _, _, 0, _, _, _, 0, 0, _, _, _, _, _, _, _,
  0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, 0, _, 0, _, _, 0, _, _, _, 0, 0, _, _, _, _, _, _, _,
  0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, 0, _, 0, _, _, 0, _, _, _, 0, 0, _, _, _, _, _, _, _,
  0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, 0, _, 0, _, _, 0, _, _, _, 0, 0, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, 0, _, 0, _, _, 0, _, _, _, 0, 0, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, 0, _, 0, _, _, 0, _, _, _, 0, 0, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, 0, _, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, 0, _, 0, _, _, 0, _, _, _, 0, 0, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, 0, _, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, 0, _, 0, _, _, 0, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, 0, _, 0, _, _, 0, _, _, _, 0, 0, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, 0, _, 0, _, _, 0, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, 0, _, 0, _, _, 0, _, _, _, 0, 0, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, 0, _, 0, _, _, 0, _, _, _, 0, 0, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, 0, _, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 Silicate =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 2.04, 1.09, 2.37, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _,
  4.201456, 4.201456, 4.196061, 4.186676, 4.165851, 4.180905, 4.201456, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4.201456, 4.201456, 4.196061, 4.186676, 4.165851, 4.180905, 4.201456, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4.201456, 4.201456, 4.196061, 4.186676, 4.165851, 4.180905, 4.201456, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4.201456, 4.201456, 4.196061, 4.186676, 4.165851, 4.180905, 4.201456, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4.201456, 4.201456, 4.196061, 4.186676, 4.165851, 4.180905, 4.201456, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4.201456, 4.201456, 4.196061, 4.186676, 4.165851, 4.180905, 4.201456, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  29.6904, 31.86794, 33.41051, 34.04187, 34.57068, 34.80565, _, _, _, _, 
    46.74787, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  29.6904, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _,
  1.6, 2.8, 1.8, 3.2, 2.8, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _,
  1.6, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  1.6, 2.8, 1.8, 3.2, 2.8, 34.80565, _, _, _, _, 46.74787, _, _, _, _, _, _, 
    112.5246, 121.2695, 129.5414, _, _, _, _, _, _,
  3.916, 7.191199, 9.967999, 11.96531, 15.308, 22.83477, 29.904, _, 42.48267, 
    53.044, _, _, _, 81.88, _, _, 97.89999, 104.7125, 112.14, 119.9275, 
    128.16, _, _, _, _, _,
  3.916, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  3.916, 7.191199, 9.967999, 11.96531, 15.308, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _,
  3.916, 7.191199, 9.967999, 11.96531, 15.308, 22.83477, 29.904, _, 42.48267, 
    53.044, _, _, _, 81.88, _, _, 97.89999, 104.7125, 112.14, 119.9275, 
    128.16, _, _, _, _, 16.03816,
  3.916, 7.191199, 9.967999, 11.96531, 15.308, 22.83477, 29.904, _, 42.48267, 
    53.044, _, _, _, 81.88, _, _, _, _, _, _, _, _, _, _, _, _,
  3.916, 7.191199, 9.967999, 11.96531, 15.308, 22.83477, 29.904, _, 42.48267, 
    53.044, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3.916, 7.191199, 9.967999, 11.96531, 15.308, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _,
  3.916, 7.191199, 9.967999, 11.96531, 15.308, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _,
  3.916, 7.191199, 9.967999, 11.96531, 15.308, 22.83477, 29.904, _, 42.48267, 
    53.044, _, _, _, 81.88, _, _, 97.89999, 104.7125, 112.14, 119.9275, 
    128.16, _, _, _, _, _,
  3.916, 7.191199, 9.967999, 11.96531, 15.308, 22.83477, 29.904, _, 42.48267, 
    53.044, _, _, _, 81.88, _, _, _, _, _, _, _, _, _, _, _, _,
  3.916, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  1.1, 2.7, 2.3, 2.2, 2.2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _,
  1.1, 2.7, 2.3, 2.2, 2.2, 22.83477, 29.904, _, 42.48267, 53.044, _, _, _, 
    81.88, _, _, 97.89999, 104.7125, 112.14, 119.9275, 128.16, _, _, _, _, _,
  1.1, 2.5, 1.6, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _,
  1.1, 2.5, 1.6, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _,
  1.1, 2.5, 1.6, 3, 2.2, 22.83477, 29.904, _, 42.48267, 53.044, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _,
  1.1, 2.5, 1.6, 3, 2.2, 22.83477, 29.904, _, 42.48267, 53.044, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _,
  1.1, 2.5, 1.6, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _,
  4, 3.9, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  4, 3.9, 1.6, 3, 2.2, 22.83477, 29.904, _, 42.48267, 53.044, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _,
  4, 3.9, 1.6, 3, 2.2, 22.83477, 29.904, _, 42.48267, 53.044, _, _, _, 81.88, 
    _, _, 97.89999, 104.7125, 112.14, 119.9275, _, _, _, _, _, _,
  8.971, 8.971, 8.971, 8.971, 8.971, 8.971, 8.971, 8.971, 8.971, 8.971, 
    8.971, 8.971, 9.968, 11.997, 12.994, 12.994, 11.997, 10.98552, 9.968, 
    11.06349, 11.997, 12.56407, 12.85674, 12.994, _, 12.994,
  8.971, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  8.971, 8.971, 8.971, 8.971, 8.971, 8.971, 8.971, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _,
  8.971, 8.971, 8.971, 8.971, 8.971, 8.971, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _,
  8.971, 8.971, 8.971, 8.971, 8.971, 8.971, 8.971, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _,
  8.971, 8.971, 8.971, 8.971, 8.971, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _,
  8.971, 8.971, 8.971, 8.971, 8.971, 8.971, 8.971, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _,
  8.971, 8.971, 8.971, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _,
  8.971, 8.971, 8.971, 8.971, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _,
  8.971, 8.971, 8.971, 8.971, 8.971, 8.971, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _,
  8.971, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  8.971, 8.971, 8.971, 8.971, 8.971, 8.971, 8.971, 8.971, 8.971, 8.971, 
    8.971, 8.971, 9.968, 11.997, 12.994, 12.994, 11.997, 10.98552, 9.968, 
    11.06349, 11.997, 12.56407, 12.85674, 12.994, _, _,
  8.971, 8.971, 8.971, 8.971, 8.971, 8.971, 8.971, 8.971, 8.971, 8.971, 
    8.971, 8.971, 9.968, 11.997, 12.994, _, _, _, _, _, _, _, _, _, _, _,
  8.971, 8.971, 8.971, 8.971, 8.971, 8.971, 8.971, 8.971, 8.971, 8.971, 
    8.971, 8.971, 9.968, 11.997, 12.994, 12.994, 11.997, 10.98552, 9.968, 
    11.06349, 11.997, _, _, _, _, _,
  5, 4.4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  5, 4.4, 8.971, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _,
  5, 4.4, 8.971, 8.971, 8.971, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _,
  5, 4.4, 8.971, 8.971, 8.971, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _,
  5, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  5, 4.4, 8.971, 8.971, 8.971, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _,
  5, 4.4, 8.971, 8.971, 8.971, 8.971, 8.971, 8.971, 8.971, 8.971, 8.971, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  5, 4.4, 8.971, 8.971, 8.971, 8.971, 8.971, 8.971, 8.971, 8.971, 8.971, 
    8.971, 9.968, 11.997, 12.994, 12.994, 11.997, 10.98552, 9.968, 11.06349, 
    11.997, 12.56407, 12.85674, 12.994, _, _,
  5, 4.4, 8.971, 8.971, 8.971, 8.971, 8.971, 8.971, 8.971, 8.971, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _,
  5, 4.4, 8.971, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _,
  4.7, 4.3, 4.7, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _,
  4.2, 4.6, 4.2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _,
  13.88617, 13.61362, 13.71662, 13.63185, 13.85677, 14.90856, 15.89812, 
    16.80818, 17.50509, 18.8579, _, _, _, _, _, _, _, _, 96.78901, _, _, _, 
    _, _, _, _,
  13.88617, 13.61362, 13.71662, 13.63185, 13.85677, 14.90856, 15.89812, 
    16.80818, 17.50509, 18.8579, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  13.88617, 13.61362, 13.71662, 13.63185, 13.85677, 14.90856, 15.89812, 
    16.80818, 17.50509, 18.8579, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  13.88617, 13.61362, 13.71662, 13.63185, 13.85677, 14.90856, 15.89812, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  13.88617, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _,
  13.88617, 13.61362, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _,
  13.88617, 13.61362, 13.71662, 13.63185, 13.85677, 14.90856, 15.89812, 
    16.80818, 17.50509, 18.8579, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4.6, 4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  4.6, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  4.6, 4, 13.71662, 13.63185, 13.85677, 14.90856, 15.89812, 16.80818, 
    17.50509, 18.8579, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4.7, 4.1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  4.7, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  4.7, 4.1, 13.71662, 13.63185, 13.85677, 14.90856, 15.89812, 16.80818, 
    17.50509, 18.8579, _, _, _, _, _, _, _, _, 96.78901, _, _, _, _, _, _, _,
  4.7, 4.1, 13.71662, 13.63185, 13.85677, 14.90856, 15.89812, 16.80818, 
    17.50509, 18.8579, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4.7, 4.1, 13.71662, 13.63185, 13.85677, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _,
  4.7, 4.1, 13.71662, 13.63185, 13.85677, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _,
  4.7, 4.1, 13.71662, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _,
  2.9, 0.9, 2.1, 1.6, 2.3, 1.7, 2.9, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _,
  2.9, 0.9, 2.1, 1.6, 2.3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _,
  2.9, 0.9, 2.1, 1.6, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _,
  3.6, 3.7, 3.633333, 3.65, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _,
  3.6, 3.7, 3.633333, 3.65, _, 1.7, 2.9, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _,
  3.6, 3.7, 3.633333, 3.65, _, 1.7, 2.9, 16.80818, 17.50509, 18.8579, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3.6, 3.7, 3.633333, 3.65, _, 1.7, 2.9, 16.80818, 17.50509, 18.8579, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  10.965, 9.968, 9.968, 10.965, 9.968, 10.965, 9.968, 11.18293, 11.997, 
    11.997, 12.994, 12.994, 12.994, 12.994, 10.965, 12.994, 13.991, 12.36042, 
    10.965, 11.05069, 11.997, 13.2964, 15.42524, 16.981, _, 16.03816,
  5.696, 10.34773, 14.24, 16.5118, 21.36, 28.35757, 35.956, _, 46.636, 53.4, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  5.696, 10.34773, 14.24, 16.5118, 21.36, 28.35757, 35.956, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _,
  5.696, 10.34773, 14.24, 16.5118, 21.36, 28.35757, 35.956, _, 46.636, 53.4, 
    12.994, 12.994, 12.994, 12.994, _, _, _, _, _, _, _, _, _, _, _, _,
  5.696, 10.34773, 14.24, 16.5118, 21.36, 28.35757, 35.956, _, 46.636, 53.4, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2.7, 3.6, 3.1, 2.6, 2.7, 2.3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _,
  2.7, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  2.7, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  2.7, 3.6, 3.1, 2.6, 2.7, 2.3, _, _, 46.636, 53.4, 12.994, 12.994, 12.994, 
    12.994, 10.965, 12.994, 13.991, 12.36042, 10.965, 11.05069, 11.997, 
    13.2964, 15.42524, 16.981, _, _,
  2.7, 3.6, 3.1, 2.6, 2.7, 2.3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _,
  2.7, 3.6, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  2.7, 3.6, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  2.7, 3.6, 3.1, 2.6, 2.7, 2.3, _, _, 46.636, 53.4, 12.994, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _,
  2.7, 3.6, 3.1, 2.6, 2.7, 2.3, _, _, 46.636, 53.4, 12.994, 12.994, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _,
  2.7, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  2.7, 3.6, 3.1, 2.6, 2.7, 2.3, _, _, 46.636, 53.4, 12.994, 12.994, 12.994, 
    12.994, 10.965, 12.994, 13.991, 12.36042, 10.965, 11.05069, 11.997, 
    13.2964, 15.42524, 16.981, _, _,
  2.7, 3.6, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  2.7, 3.6, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  2.7, 3.6, 3.1, 2.6, 2.7, 2.3, _, _, 46.636, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _,
  2.7, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  2.7, 3.6, 3.1, 2.6, 2.7, 2.3, _, _, 46.636, 53.4, 12.994, 12.994, 12.994, 
    12.994, 10.965, 12.994, 13.991, 12.36042, 10.965, 11.05069, 11.997, 
    13.2964, 15.42524, 16.981, _, _,
  2.7, 3.6, 3.1, 2.6, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _,
  2.7, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  2.7, 3.6, 3.1, 2.6, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _,
  2.7, 3.6, 3.1, 2.6, 2.7, 2.3, _, _, 46.636, 53.4, 12.994, 12.994, 12.994, 
    12.994, 10.965, 12.994, 13.991, 12.36042, 10.965, 11.05069, 11.997, 
    13.2964, 15.42524, 16.981, _, 16.03816,
  2.7, 3.6, 3.1, 2.6, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _,
  2.7, 3.6, 3.1, 2.6, 2.7, 2.3, _, _, 46.636, 53.4, 12.994, 12.994, 12.994, 
    12.994, 10.965, 12.994, 13.991, 12.36042, 10.965, 11.05069, _, _, _, _, 
    _, _,
  2.7, 3.6, 3.1, 2.6, 2.7, 2.3, _, _, 46.636, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _,
  2.7, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  2.7, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  2.7, 3.6, 3.1, 2.6, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _,
  2.7, 3.6, 3.1, 2.6, 2.7, 2.3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _,
  2.7, 3.6, 3.1, 2.6, 2.7, 2.3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _,
  2.7, 3.6, 3.1, 2.6, 2.7, 2.3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _,
  2.7, 3.6, 3.1, 2.6, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _,
  2.7, 3.6, 3.1, 2.6, 2.7, 2.3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _,
  2.7, 3.6, 3.1, 2.6, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _,
  2.7, 3.6, 3.1, 2.6, 2.7, 2.3, _, _, 46.636, 53.4, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _,
  11.74984, 12.06174, 12.38481, 12.71903, 13.42097, 14.36307, 15.41747, 
    16.22099, 16.8588, 17.65024, 18.05427, _, _, _, _, _, _, _, 98.99327, 
    105.5264, _, _, _, _, _, _,
  8.9, 14.00267, 18.156, 20.97476, 24.92, 37.38, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _,
  8.9, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  8.9, 14.00267, 18.156, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _,
  8.9, 14.00267, 18.156, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _,
  8.9, 14.00267, 18.156, 20.97476, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _,
  8.9, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  8.9, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  8.9, 14.00267, 18.156, 20.97476, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _,
  8.9, 14.00267, 18.156, 20.97476, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _,
  8.9, 14.00267, 18.156, 20.97476, 24.92, 37.38, 15.41747, 16.22099, 16.8588, 
    17.65024, 18.05427, _, _, _, _, _, _, _, 98.99327, 105.5264, _, _, _, _, 
    _, _,
  8.9, 14.00267, 18.156, 20.97476, 24.92, 37.38, 15.41747, 16.22099, 16.8588, 
    17.65024, 18.05427, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  8.9, 14.00267, 18.156, 20.97476, 24.92, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _,
  8.9, 14.00267, 18.156, 20.97476, 24.92, 37.38, 15.41747, 16.22099, 16.8588, 
    17.65024, 18.05427, _, _, _, _, _, _, _, 98.99327, 105.5264, _, _, _, _, 
    _, _,
  8.9, 14.00267, 18.156, 20.97476, 24.92, 37.38, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _,
  8.9, 14.00267, 18.156, 20.97476, 24.92, 37.38, 15.41747, 16.22099, 16.8588, 
    17.65024, 18.05427, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  8.9, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  8.9, 14.00267, 18.156, 20.97476, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _,
  8.9, 14.00267, 18.156, 20.97476, 24.92, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _,
  8.9, 14.00267, 18.156, 20.97476, 24.92, 37.38, 15.41747, 16.22099, 16.8588, 
    17.65024, 18.05427, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  8.9, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  8.9, 14.00267, 18.156, 20.97476, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _,
  8.9, 14.00267, 18.156, 20.97476, 24.92, 37.38, 15.41747, 16.22099, 16.8588, 
    17.65024, 18.05427, _, _, _, _, _, _, _, 98.99327, 105.5264, _, _, _, _, 
    _, _,
  8.9, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  8.9, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  8.9, 14.00267, 18.156, 20.97476, 24.92, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _,
  8.9, 14.00267, 18.156, 20.97476, 24.92, 37.38, 15.41747, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _,
  8.9, 14.00267, 18.156, 20.97476, 24.92, 37.38, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _,
  8.9, 14.00267, 18.156, 20.97476, 24.92, 37.38, 15.41747, 16.22099, 16.8588, 
    17.65024, 18.05427, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4.272, 9.885791, 14.22835, 16.05466, 20.74993, 29.09345, _, _, _, _, _, _, 
    _, _, _, _, _, 112.5246, 121.2695, 129.5414, _, _, _, _, _, _,
  4.272, 9.885791, 14.22835, 16.05466, 20.74993, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _,
  4.272, 9.885791, 14.22835, 16.05466, 20.74993, 29.09345, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4.272, 9.885791, 14.22835, 16.05466, 20.74993, 29.09345, _, _, _, _, _, _, 
    _, _, _, _, _, 112.5246, 121.2695, 129.5414, _, _, _, _, _, _,
  3.9, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  5.1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  2.7, 2.5, 2.7, 2.2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _,
  5.5, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  5.5, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  3.3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  3.3, 2.5, 2.7, 2.2, 20.74993, 29.09345, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _,
  3.4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  4.8, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  3.6, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  3.3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _ ;

 Silicate_sigfigs =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 4, 4, 4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  5, 5, 5, 5, 5, 5, 5, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  5, 5, 5, 5, 5, 5, 5, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  5, 5, 5, 5, 5, 5, 5, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  5, 5, 5, 5, 5, 5, 5, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  5, 5, 5, 5, 5, 5, 5, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  5, 5, 5, 5, 5, 5, 5, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 3, 3, 3, 3, 3, _, _, _, _, 4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, 2, 3, _, _, _, _, 4, _, _, _, _, _, _, 5, 5, 5, _, _, _, _, _, _,
  1, 4, 4, 4, 4, 4, 4, _, 4, 5, _, _, _, 5, _, _, 5, 5, 5, 5, 5, _, _, _, _, _,
  1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, 4, 4, 4, 4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, 4, 4, 4, 4, 4, 4, _, 4, 5, _, _, _, 5, _, _, 5, 5, 5, 5, 5, _, _, _, _, 5,
  1, 4, 4, 4, 4, 4, 4, _, 4, 5, _, _, _, 5, _, _, _, _, _, _, _, _, _, _, _, _,
  1, 4, 4, 4, 4, 4, 4, _, 4, 5, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, 4, 4, 4, 4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, 4, 4, 4, 4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, 4, 4, 4, 4, 4, 4, _, 4, 5, _, _, _, 5, _, _, 5, 5, 5, 5, 5, _, _, _, _, _,
  1, 4, 4, 4, 4, 4, 4, _, 4, 5, _, _, _, 5, _, _, _, _, _, _, _, _, _, _, _, _,
  1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, 2, 4, 4, _, 4, 5, _, _, _, 5, _, _, 5, 5, 5, 5, 5, _, _, _, _, _,
  2, 2, 2, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, 2, 4, 4, _, 4, 5, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, 2, 4, 4, _, 4, 5, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, 2, 4, 4, _, 4, 5, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, 2, 4, 4, _, 4, 5, _, _, _, 5, _, _, 5, 5, 5, 5, _, _, _, _, _, _,
  4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 5, 5, 5, 5, 5, 4, 5, 5, 5, 5, 5, _, 5,
  4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4, 4, 4, 4, 4, 4, 4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4, 4, 4, 4, 4, 4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4, 4, 4, 4, 4, 4, 4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4, 4, 4, 4, 4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4, 4, 4, 4, 4, 4, 4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4, 4, 4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4, 4, 4, 4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4, 4, 4, 4, 4, 4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 5, 5, 5, 5, 5, 4, 5, 5, 5, 5, 5, _, _,
  4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 5, 5, _, _, _, _, _, _, _, _, _, _, _,
  4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 5, 5, 5, 5, 5, 4, 5, 5, _, _, _, _, _,
  2, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 4, 4, 4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 4, 4, 4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 4, 4, 4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 4, 4, 4, 4, 4, 4, 4, 4, 4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 5, 5, 5, 5, 5, 4, 5, 5, 5, 5, 5, _, _,
  2, 2, 4, 4, 4, 4, 4, 4, 4, 4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 4, 4, 4, 4, 4, 4, 4, 4, 4, _, _, _, _, _, _, _, _, 4, _, _, _, _, _, _, _,
  2, 4, 4, 4, 4, 4, 4, 4, 4, 4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 4, 4, 4, 4, 4, 4, 4, 4, 4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 4, 4, 4, 4, 4, 4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 4, 4, 4, 4, 4, 4, 4, 4, 4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 4, 4, 4, 4, 4, 4, 4, 4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 4, 4, 4, 4, 4, 4, 4, 4, _, _, _, _, _, _, _, _, 4, _, _, _, _, _, _, _,
  2, 2, 4, 4, 4, 4, 4, 4, 4, 4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 4, 4, 4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 4, 4, 4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 1, 2, 2, 2, 2, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 1, 2, 2, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 1, 2, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, _, 2, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, _, 2, 2, 4, 4, 4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, _, 2, 2, 4, 4, 4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  5, 4, 4, 5, 4, 5, 4, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, _, 5,
  1, 4, 4, 4, 4, 4, 5, _, 5, 5, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, 4, 4, 4, 4, 4, 5, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, 4, 4, 4, 4, 4, 5, _, 5, 5, 5, 5, 5, 5, _, _, _, _, _, _, _, _, _, _, _, _,
  1, 4, 4, 4, 4, 4, 5, _, 5, 5, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, 2, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, 2, 2, _, _, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, _, _,
  2, 2, 2, 2, 2, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, 2, 2, _, _, 5, 5, 5, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, 2, 2, _, _, 5, 5, 5, 5, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, 2, 2, _, _, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, _, _,
  2, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, 2, 2, _, _, 5, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, 2, 2, _, _, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, _, _,
  2, 2, 2, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, 2, 2, _, _, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, _, 5,
  2, 2, 2, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, 2, 2, _, _, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, _, _, _, _, _, _,
  2, 2, 2, 2, 2, 2, _, _, 5, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, 2, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, 2, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, 2, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, 2, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, 2, 2, _, _, 5, 5, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, _, _, _, _, _, _, _, 4, 5, _, _, _, _, _, _,
  1, 4, 4, 4, 4, 5, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, 4, 4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, 4, 4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, 4, 4, 4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, 4, 4, 4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, 4, 4, 4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, 4, 4, 4, 4, 5, 4, 4, 4, 4, 4, _, _, _, _, _, _, _, 4, 5, _, _, _, _, _, _,
  1, 4, 4, 4, 4, 5, 4, 4, 4, 4, 4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, 4, 4, 4, 4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, 4, 4, 4, 4, 5, 4, 4, 4, 4, 4, _, _, _, _, _, _, _, 4, 5, _, _, _, _, _, _,
  1, 4, 4, 4, 4, 5, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, 4, 4, 4, 4, 5, 4, 4, 4, 4, 4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, 4, 4, 4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, 4, 4, 4, 4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, 4, 4, 4, 4, 5, 4, 4, 4, 4, 4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, 4, 4, 4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, 4, 4, 4, 4, 5, 4, 4, 4, 4, 4, _, _, _, _, _, _, _, 4, 5, _, _, _, _, _, _,
  1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, 4, 4, 4, 4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, 4, 4, 4, 4, 5, 4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, 4, 4, 4, 4, 5, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, 4, 4, 4, 4, 5, 4, 4, 4, 4, 4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, 3, 4, 4, 4, 4, _, _, _, _, _, _, _, _, _, _, _, 5, 5, 5, _, _, _, _, _, _,
  1, 3, 4, 4, 4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, 3, 4, 4, 4, 4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, 3, 4, 4, 4, 4, _, _, _, _, _, _, _, _, _, _, _, 5, 5, 5, _, _, _, _, _, _,
  1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, 4, 4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 Silicate_WODflag =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, _, _, _, _, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, _, _, _, _, 0, _, _, _, _, _, _, 0, 0, 0, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, 0, 0, _, _, _, 0, _, _, 0, 0, 0, 0, 0, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, 0, 0, _, _, _, 0, _, _, 0, 0, 0, 0, 0, _, _, _, _, 0,
  0, 0, 0, 0, 0, 0, 0, _, 0, 0, _, _, _, 0, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, 0, 0, _, _, _, 0, _, _, 0, 0, 0, 0, 0, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, 0, 0, _, _, _, 0, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, 0, 0, _, _, _, 0, _, _, 0, 0, 0, 0, 0, _, _, _, _, _,
  0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, 0, 0, _, _, _, 0, _, _, 0, 0, 0, 0, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, 0,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _,
  0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  6, 6, 6, 6, 6, 6, 6, 6, 6, 6, _, _, _, _, _, _, _, _, 6, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, 0, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, _, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, _, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, _, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, _, 0,
  0, 0, 0, 0, 0, 0, 0, _, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, _, _, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _,
  0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, _, _, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, _, _, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, _, _, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _,
  0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, _, _, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, _, _, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _,
  0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, _, _, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, 0,
  0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, _, _, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, _, _, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, _, _, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, _, _, _, _, _, _, _, 0, 6, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, 0, 0, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, 0, 0, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, 0, 0, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, 0, 0, 0, _, _, _, _, _, _,
  0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, 0, 0, 0, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 Silicate_WODprofileflag = _, _, _, _, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0 ;

 Silicate_Original_units =
  "\"ug/l\"    Alternate Nutrient Conversion (use instead of #36)",
  "\"ug/l\"    Alternate Nutrient Conversion (use instead of #36)",
  "ug/l               mg/m3    ppb     g/1000m3",
  "\"ug/l\"    Alternate Nutrient Conversion (use instead of #36)",
  "ug/l               mg/m3    ppb     g/1000m3",
  "\"ug/l\"    Alternate Nutrient Conversion (use instead of #36)",
  "ug/l               mg/m3    ppb     g/1000m3",
  "ug/l               mg/m3    ppb     g/1000m3",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "" ;

 Nitrite =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0.2141832, 0.1427888, 0.1427888, 0.1427888, 0.1427888, 0.1427888, 
    0.1427888, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0.2141832, 0.1427888, 0.1427888, 0.1427888, 0.1427888, 0.1427888, 
    0.1427888, 0.004844075, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  0.2141832, 0.1427888, 0.1427888, 0.1427888, 0.1427888, 0.1427888, 
    0.1427888, 0.004844075, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  0.2141832, 0.1427888, 0.1427888, 0.1427888, 0.1427888, 0.1427888, 
    0.1427888, 0.004844075, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  0.2141832, 0.1427888, 0.1427888, 0.1427888, 0.1427888, 0.1427888, 
    0.1427888, 0.004844075, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  0.2141832, 0.1427888, 0.1427888, 0.1427888, 0.1427888, 0.1427888, 
    0.1427888, 0.004844075, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  0.2141832, 0.1427888, 0.1427888, 0.1427888, 0.1427888, 0.1427888, 
    0.1427888, 0.004844075, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  0.2141832, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _,
  0.2141832, 0.1427888, 0.1427888, 0.1427888, 0.1427888, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0.2141832, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _,
  0.2141832, 0.1427888, 0.1427888, 0.1427888, 0.1427888, 0.1427888, 
    0.1427888, 0.004844075, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  0.2141832, 0.1427888, 0.1427888, 0.1427888, 0.1427888, 0.1427888, 
    0.1427888, 0.004844075, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  0.2141832, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _,
  0.2141832, 0.1427888, 0.1427888, 0.1427888, 0.1427888, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0.2141832, 0.1427888, 0.1427888, 0.1427888, 0.1427888, 0.1427888, 
    0.1427888, 0.004844075, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  0.2141832, 0.1427888, 0.1427888, 0.1427888, 0.1427888, 0.1427888, 
    0.1427888, 0.004844075, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  0.2141832, 0.1427888, 0.1427888, 0.1427888, 0.1427888, 0.1427888, 
    0.1427888, 0.004844075, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  0.2141832, 0.1427888, 0.1427888, 0.1427888, 0.1427888, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0.2141832, 0.1427888, 0.1427888, 0.1427888, 0.1427888, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0.2141832, 0.1427888, 0.1427888, 0.1427888, 0.1427888, 0.1427888, 
    0.1427888, 0.004844075, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  0.2141832, 0.1427888, 0.1427888, 0.1427888, 0.1427888, 0.1427888, 
    0.1427888, 0.004844075, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  0.2141832, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _,
  0.2141832, 0.1427888, 0.1427888, 0.1427888, 0.1427888, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0.2141832, 0.1427888, 0.1427888, 0.1427888, 0.1427888, 0.1427888, 
    0.1427888, 0.004844075, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  0.2141832, 0.1427888, 0.1427888, 0.1427888, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _,
  0.2141832, 0.1427888, 0.1427888, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _,
  0.2141832, 0.1427888, 0.1427888, 0.1427888, 0.1427888, 0.1427888, 
    0.1427888, 0.004844075, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  0.2141832, 0.1427888, 0.1427888, 0.1427888, 0.1427888, 0.1427888, 
    0.1427888, 0.004844075, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  0.2141832, 0.1427888, 0.1427888, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _,
  0.2141832, 0.1427888, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _,
  0.2141832, 0.1427888, 0.1427888, 0.1427888, 0.1427888, 0.1427888, 
    0.1427888, 0.004844075, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  0.2141832, 0.1427888, 0.1427888, 0.1427888, 0.1427888, 0.1427888, 
    0.1427888, 0.004844075, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  0.2141832, 0.1427888, 0.1427888, 0.1427888, 0.1427888, 0.1427888, 
    0.1427888, 0.004844075, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  0.2141832, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _,
  0.2141832, 0.1427888, 0.1427888, 0.1427888, 0.1427888, 0.1427888, 
    0.1427888, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0.2141832, 0.1427888, 0.1427888, 0.1427888, 0.1427888, 0.1427888, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0.26, 0.24, 0.19, 0.12, 0.09, 0.07017858, 0.07, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _,
  0.26, 0.24, 0.19, 0.12, 0.09, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _,
  0.26, 0.24, 0.19, 0.12, 0.09, 0.07017858, 0.07, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _,
  0.26, 0.24, 0.19, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _,
  0.26, 0.24, 0.19, 0.12, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _,
  0.07, 0.32, 0.2, 0.17, 0.07, 0.09, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _,
  0.07, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  0.07, 0.32, 0.2, 0.17, 0.07, 0.09, 0.07, 0.004844075, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _,
  0.07, 0.32, 0.2, 0.17, 0.07, 0.09, 0.07, 0.004844075, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _,
  0.07, 0.32, 0.2, 0.17, 0.07, 0.09, 0.07, 0.004844075, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _,
  0.07, 0.32, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _,
  0.07, 0.32, 0.2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _,
  0.07, 0.32, 0.2, 0.17, 0.07, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _,
  0.07, 0.32, 0.2, 0.17, 0.07, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _,
  0.07, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  0.07, 0.32, 0.2, 0.17, 0.07, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _,
  0.07, 0.32, 0.2, 0.17, 0.07, 0.09, 0.07, 0.004844075, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _,
  0.07, 0.32, 0.2, 0.17, 0.07, 0.09, 0.07, 0.004844075, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _,
  0.24, 0.19, 0.32, 0.12, 0.1, 0.07896552, 0.07, 0.08121951, 0.09, 0.07, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0.24, 0.19, 0.32, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _,
  0.24, 0.19, 0.32, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _,
  0.24, 0.19, 0.32, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _,
  0.24, 0.19, 0.32, 0.12, 0.1, 0.07896552, 0.07, 0.08121951, 0.09, 0.07, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0.24, 0.19, 0.32, 0.12, 0.1, 0.07896552, 0.07, 0.08121951, 0.09, 0.07, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0.17, 0.36, 0.17, 0.09, 0.05, 0.05, 0.05, 0.1139706, 0.2, 0.1, _, 
    0.09473684, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0.17, 0.36, 0.17, 0.09, 0.05, 0.05, 0.05, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _,
  0.17, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  0.17, 0.36, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _,
  0.17, 0.36, 0.17, 0.09, 0.05, 0.05, 0.05, 0.1139706, 0.2, 0.1, _, 
    0.09473684, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0.17, 0.36, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _,
  0.17, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  0.37, 0.14, 0.15, 0.09, 0.12, 0.09270638, 0.07, 0.06, 0.05, 0.03, _, 
    0.03200001, 0.09, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0.37, 0.14, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _,
  0.37, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  0.37, 0.14, 0.15, 0.09, 0.12, 0.09270638, 0.07, 0.06, 0.05, 0.03, _, 
    0.03200001, 0.09, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0.37, 0.14, 0.15, 0.09, 0.12, 0.09270638, 0.07, 0.06, 0.05, 0.03, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _,
  0.37, 0.14, 0.15, 0.09, 0.12, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _,
  0.37, 0.14, 0.15, 0.09, 0.12, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _,
  0.03, _, 0.02363636, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _,
  0.03, _, 0.02363636, 0.09, 0.12, 0.09270638, 0.07, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _,
  0.03, _, 0.02363636, 0.09, 0.12, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _,
  0.03, _, 0.02363636, 0.09, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _,
  0.03, _, 0.02363636, 0.09, 0.12, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _,
  0.03, _, 0.02363636, 0.09, 0.12, 0.09270638, 0.07, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _,
  0.1, 0.12, 0.14, 0.17, 0.09, 0.09569575, 0.1, 0.09827273, 0.09, 0.05, _, 
    0.08499999, 0.12, 0.11, 0.07, _, _, _, _, _, _, _, _, _, _, _,
  0.1, 0.12, 0.14, 0.17, 0.09, 0.09569575, 0.1, 0.09827273, 0.09, 0.05, _, 
    0.08499999, 0.12, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0.1, 0.12, 0.14, 0.17, 0.09, 0.09569575, 0.1, 0.09827273, 0.09, 0.05, _, 
    0.08499999, 0.12, 0.11, 0.07, _, _, _, _, _, _, _, _, _, _, _,
  0.1, 0.12, 0.14, 0.17, 0.09, 0.09569575, 0.1, 0.09827273, 0.09, 0.05, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0.1, 0.12, 0.14, 0.17, 0.09, 0.09569575, 0.1, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _,
  0.1, 0.12, 0.14, 0.17, 0.09, 0.09569575, 0.1, 0.09827273, 0.09, 0.05, _, 
    0.08499999, 0.12, 0.11, _, _, _, _, _, _, _, _, _, _, _, _,
  0.1, 0.12, 0.14, 0.17, 0.09, 0.09569575, 0.1, 0.09827273, 0.09, 0.05, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0.1, 0.12, 0.14, 0.17, 0.09, 0.09569575, 0.1, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _,
  0.1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  0.1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  0.1, 0.12, 0.14, 0.17, 0.09, 0.09569575, 0.1, 0.09827273, 0.09, 0.05, _, 
    0.08499999, 0.12, 0.11, 0.07, _, _, _, _, _, _, _, _, _, _, _,
  0.1, 0.12, 0.14, 0.17, 0.09, 0.09569575, 0.1, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _,
  0.1, 0.12, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _,
  0.1, 0.12, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _,
  0.1, 0.12, 0.14, 0.17, 0.09, 0.09569575, 0.1, 0.09827273, 0.09, 0.05, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0.1, 0.29, 0.63, 0.24, 0.17, 0.1602459, 0.15, 0.1351793, 0.12, 0.34, _, 
    0.2136842, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0.1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  0.1, 0.29, 0.63, 0.24, 0.17, 0.1602459, 0.15, 0.1351793, 0.12, 0.34, _, 
    0.2136842, 0.12, 0.11, 0.07, _, _, _, _, _, _, _, _, _, _, _,
  0.1, 0.29, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _,
  0.1, 0.29, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _,
  0.1, 0.29, 0.63, 0.24, 0.17, 0.1602459, 0.15, 0.1351793, 0.12, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _,
  0.1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  0.1, 0.29, 0.63, 0.24, 0.17, 0.1602459, 0.15, 0.1351793, 0.12, 0.34, _, 
    0.2136842, 0.12, 0.11, 0.07, _, _, _, _, _, _, _, _, _, _, _,
  0.02, 0.002, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _,
  0.02, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  0.02, 0.002, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _,
  0.02, 0.002, _, _, 0.17, 0.1602459, 0.15, 0.1351793, 0.12, 0.34, _, 
    0.2136842, 0.12, 0.11, 0.07, _, _, _, _, _, _, _, _, _, _, _,
  0.02, 0.002, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _,
  0.02, 0.002, _, _, 0.17, 0.1602459, 0.15, 0.1351793, 0.12, 0.34, _, 
    0.2136842, 0.12, 0.11, 0.07, _, _, _, _, _, _, _, _, _, _, _,
  0.07, 0.29, 0.09, 0.09, 0.07, 0.07, 0.07, 0.085, 0.1, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _,
  0.07, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  0.07, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  0.07, 0.29, 0.09, 0.09, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _,
  _, _, _, _, 0.1172573, 0.18, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _,
  _, _, _, _, 0.1172573, 0.18, 0.07, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _,
  0.17, 0.46, 0.24, 0.1, 0.07, 0.08071429, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _,
  0.17, 0.46, 0.24, 0.1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _,
  0.17, 0.46, 0.24, 0.1, 0.07, 0.08071429, 0.07, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _,
  0.17, 0.46, 0.24, 0.1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _,
  0.17, 0.46, 0.24, 0.1, 0.07, 0.08071429, 0.07, 0.085, 0.1, 0.34, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _,
  0.17, 0.46, 0.24, 0.1, 0.07, 0.08071429, 0.07, 0.085, 0.1, 0.34, _, 
    0.2136842, 0.12, 0.11, 0.07, _, _, _, _, _, _, _, _, _, _, _,
  0.17, 0.46, 0.24, 0.1, 0.07, 0.08071429, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _,
  0.17, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  0.17, 0.46, 0.24, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _,
  0.17, 0.46, 0.24, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _,
  0.07, 0.2, 0.15, 0.15, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _,
  0.07, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  0.07, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  0.07, 0.2, 0.15, 0.15, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _,
  0.07, 0.2, 0.15, 0.15, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _,
  0.07, 0.2, 0.15, 0.15, 0.07, 0.08071429, 0.07, 0.085, 0.1, 0.34, _, 
    0.2136842, 0.12, 0.11, 0.07, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, 0.1285336, 0.4880708, _, 0.01622618, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _,
  1.02, 0.83, 0.7, 0.43, 0.22, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _,
  1.02, 0.83, 0.7, 0.43, 0.22, 0.4880708, _, 0.01622618, _, _, _, _, 0.12, 
    0.11, 0.07, _, _, _, _, _, _, _, _, _, _, _,
  1.02, 0.83, 0.7, 0.43, 0.22, 0.4880708, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _,
  1.02, 0.83, 0.7, 0.43, 0.22, 0.4880708, _, 0.01622618, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _,
  1.02, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  1.02, 0.83, 0.7, 0.43, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _,
  1.02, 0.83, 0.7, 0.43, 0.22, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _,
  _, _, _, _, 0.07, 0.34, 0.02, 0.004844075, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, 0.07, 0.34, 0.02, 0.004844075, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, 0.07, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  _, _, _, _, 0.07, 0.34, 0.02, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _,
  _, _, _, _, 0.07, 0.34, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _,
  _, _, _, _, 0.07, 0.34, 0.02, 0.004844075, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _,
  _, _, _, _, 0.07, 0.34, 0.02, 0.004844075, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _,
  _, _, _, _, 0.07, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  _, _, _, _, 0.07, 0.34, 0.02, 0.004844075, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _,
  _, _, _, _, 0.07, 0.34, 0.02, 0.004844075, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _,
  0.16, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  0.39, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  0.39, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  0.17, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  0.17, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  0.22, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  0.22, _, _, _, 0.07, 0.34, 0.02, 0.004844075, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _,
  0.25, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  0.17, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  0.17, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  0.22, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _ ;

 Nitrite_sigfigs =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, 3, 3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, 3, 3, 3, 3, 3, 1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, 3, 3, 3, 3, 3, 1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, 3, 3, 3, 3, 3, 1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, 3, 3, 3, 3, 3, 1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, 3, 3, 3, 3, 3, 1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, 3, 3, 3, 3, 3, 1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, 3, 3, 3, 3, 3, 1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, 3, 3, 3, 3, 3, 1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, 3, 3, 3, 3, 3, 1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, 3, 3, 3, 3, 3, 1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, 3, 3, 3, 3, 3, 1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, 3, 3, 3, 3, 3, 1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, 3, 3, 3, 3, 3, 1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, 3, 3, 3, 3, 3, 1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, 3, 3, 3, 3, 3, 1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, 3, 3, 3, 3, 3, 1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, 3, 3, 3, 3, 3, 1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, 3, 3, 3, 3, 3, 1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, 3, 3, 3, 3, 3, 1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, 3, 3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, 3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, 2, 2, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, 2, 2, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, 2, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, 2, 2, 2, 1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, 2, 2, 2, 1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, 2, 2, 2, 1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, 2, 2, 2, 1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, 2, 2, 2, 1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, 2, 2, 2, 2, 2, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, 2, 2, 2, 2, 2, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, 2, 2, 2, 2, 2, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, 2, 2, 2, 2, 2, 2, _, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, 2, 2, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, 2, 2, 2, 2, 2, 2, _, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, 2, 2, 2, 2, 2, 2, _, 2, 2, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, 2, 2, 2, 2, 2, 2, _, 2, 2, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, 2, 2, 2, 2, 2, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, _, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, _, 2, 2, 2, 2, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, _, 2, 2, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, _, 2, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, _, 2, 2, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, _, 2, 2, 2, 2, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, 2, 2, 2, 2, 2, 2, _, 2, 2, 2, 2, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, 2, 2, 2, 2, 2, 2, _, 2, 2, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, 2, 2, 2, 2, 2, 2, _, 2, 2, 2, 2, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, 2, 2, 2, 2, 2, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, 2, 2, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, 2, 2, 2, 2, 2, 2, _, 2, 2, 2, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, 2, 2, 2, 2, 2, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, 2, 2, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, 2, 2, 2, 2, 2, 2, _, 2, 2, 2, 2, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, 2, 2, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, 2, 2, 2, 2, 2, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, 2, 2, 2, 2, 2, 2, _, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, 2, 2, 2, 2, 2, 2, _, 2, 2, 2, 2, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, 2, 2, 2, 2, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, 2, 2, 2, 2, 2, 2, _, 2, 2, 2, 2, _, _, _, _, _, _, _, _, _, _, _,
  1, 1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, 1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, 1, _, _, 2, 2, 2, 2, 2, 2, _, 2, 2, 2, 2, _, _, _, _, _, _, _, _, _, _, _,
  1, 1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, 1, _, _, 2, 2, 2, 2, 2, 2, _, 2, 2, 2, 2, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, 2, 2, 2, 2, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, 2, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, 2, 2, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, 2, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, 2, 2, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, 2, 2, 2, 2, 2, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, 2, 2, 2, 2, 2, 2, _, 2, 2, 2, 2, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, 2, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, 2, 2, 2, 2, 2, 2, _, 2, 2, 2, 2, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, 1, 2, _, 1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 2, 2, 2, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 2, 2, 2, 2, 2, _, 1, _, _, _, _, 2, 2, 2, _, _, _, _, _, _, _, _, _, _, _,
  3, 2, 2, 2, 2, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 2, 2, 2, 2, 2, _, 1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 2, 2, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 2, 2, 2, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, 2, 2, 2, 1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, 2, 2, 2, 1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, 2, 2, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, 2, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, 2, 2, 2, 1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, 2, 2, 2, 1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, 2, 2, 2, 1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, 2, 2, 2, 1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, _, _, _, 2, 2, 2, 1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 Nitrite_WODflag =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, _, _, 0, 0, 0, 0, 0, 0, _, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, _, _, 0, 0, 0, 0, 0, 0, _, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, 0, 0, _, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, _, 0, _, _, _, _, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, _, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 Nitrite_Original_units =
  "\"ug/l\"    Alternate Nutrient Conversion (use instead of #36)",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "" ;

 Nitrate =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3.998087, 4.926214, 5.173376, 5.225662, 5.35458, 5.460759, 5.497369, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3.998087, 4.926214, 5.173376, 5.225662, 5.35458, 5.460759, 5.497369, 
    7.871645, 7.8, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3.998087, 4.926214, 5.173376, 5.225662, 5.35458, 5.460759, 5.497369, 
    7.871645, 7.8, 16.0435, 16.57422, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  3.998087, 4.926214, 5.173376, 5.225662, 5.35458, 5.460759, 5.497369, 
    7.871645, 7.8, 16.0435, 16.57422, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  3.998087, 4.926214, 5.173376, 5.225662, 5.35458, 5.460759, 5.497369, 
    7.871645, 7.8, 16.0435, 16.57422, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  3.998087, 4.926214, 5.173376, 5.225662, 5.35458, 5.460759, 5.497369, 
    7.871645, 7.8, 16.0435, 16.57422, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  3.998087, 4.926214, 5.173376, 5.225662, 5.35458, 5.460759, 5.497369, 
    7.871645, 7.8, 16.0435, 16.57422, 17.12065, 20.44291, _, _, _, _, _, _, 
    _, _, _, _, _, _, _,
  3.998087, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _,
  2.3, 4.4, 2.7, 3.8, 4.2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _,
  2.3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  2.3, 4.4, 2.7, 3.8, 4.2, 5.460759, 5.497369, 7.871645, 7.8, 16.0435, 
    16.57422, 17.12065, 20.44291, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2.3, 4.4, 2.7, 3.8, 4.2, 5.460759, 5.497369, 7.871645, 7.8, 16.0435, 
    16.57422, 17.12065, 20.44291, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2.3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  2.3, 4.4, 2.7, 3.8, 4.2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _,
  2.3, 4.4, 2.7, 3.8, 4.2, 5.460759, 5.497369, 7.871645, 7.8, 16.0435, 
    16.57422, 17.12065, 20.44291, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2.3, 4.4, 2.7, 3.8, 4.2, 5.460759, 5.497369, 7.871645, 7.8, 16.0435, 
    16.57422, 17.12065, 20.44291, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2.3, 4.4, 2.7, 3.8, 4.2, 5.460759, 5.497369, 7.871645, 7.8, 16.0435, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2.3, 4.4, 2.7, 3.8, 4.2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _,
  2.3, 4.4, 2.7, 3.8, 4.2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _,
  2.3, 4.4, 2.7, 3.8, 4.2, 5.460759, 5.497369, 7.871645, 7.8, 16.0435, 
    16.57422, 17.12065, 20.44291, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2.3, 4.4, 2.7, 3.8, 4.2, 5.460759, 5.497369, 7.871645, 7.8, 16.0435, 
    16.57422, 17.12065, 20.44291, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2.3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  1.9, 4.9, 3.3, 3.1, 2.7, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _,
  1.9, 4.9, 3.3, 3.1, 2.7, 5.460759, 5.497369, 7.871645, 7.8, 16.0435, 
    16.57422, 17.12065, 20.44291, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1.6, 3.2, 2.2, 3.8, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _,
  1.6, 3.2, 2.2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _,
  1.6, 3.2, 2.2, 3.8, 2.7, 5.460759, 5.497369, 7.871645, 7.8, 16.0435, 
    16.57422, 17.12065, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1.6, 3.2, 2.2, 3.8, 2.7, 5.460759, 5.497369, 7.871645, 7.8, 16.0435, 
    16.57422, 17.12065, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1.6, 3.2, 2.2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _,
  7, 7.5, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  7, 7.5, 2.2, 3.8, 2.7, 5.460759, 5.497369, 7.871645, 7.8, 16.0435, 
    16.57422, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  7, 7.5, 2.2, 3.8, 2.7, 5.460759, 5.497369, 7.871645, 7.8, 16.0435, 
    16.57422, 17.12065, 20.44291, _, _, _, _, _, _, _, _, _, _, _, _, _,
  7, 7.5, 2.2, 3.8, 2.7, 5.460759, 5.497369, 7.871645, 7.8, 16.0435, 
    16.57422, 17.12065, 20.44291, _, _, _, _, _, _, _, _, _, _, _, _, _,
  7, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  7, 7.5, 2.2, 3.8, 2.7, 5.460759, 5.497369, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _,
  7, 7.5, 2.2, 3.8, 2.7, 5.460759, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _,
  3.8, 3.8, 6.5, 8.2, 6.8, 7.45, 8.1, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _,
  3.8, 3.8, 6.5, 8.2, 6.8, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _,
  3.8, 3.8, 6.5, 8.2, 6.8, 7.45, 8.1, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _,
  3.8, 3.8, 6.5, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _,
  3.8, 3.8, 6.5, 8.2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _,
  0.3, 5.4, 7.2, 10.2, 5.9, 9.4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _,
  0.3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  0.3, 5.4, 7.2, 10.2, 5.9, 9.4, 8.1, 7.871645, 7.8, 16.0435, 16.57422, 
    17.12065, 20.44291, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0.3, 5.4, 7.2, 10.2, 5.9, 9.4, 8.1, 7.871645, 7.8, 16.0435, 16.57422, 
    17.12065, 20.44291, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0.3, 5.4, 7.2, 10.2, 5.9, 9.4, 8.1, 7.871645, 7.8, 16.0435, 16.57422, 
    17.12065, 20.44291, _, _, _, _, _, _, _, _, _, _, _, _, _,
  6, 9.4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  6, 9.4, 7.2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  6, 9.4, 7.2, 10.2, 5.9, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _,
  6, 9.4, 7.2, 10.2, 5.9, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _,
  6, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  6, 9.4, 7.2, 10.2, 5.9, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _,
  6, 9.4, 7.2, 10.2, 5.9, 9.4, 8.1, 7.871645, 7.8, 16.0435, 16.57422, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _,
  6, 9.4, 7.2, 10.2, 5.9, 9.4, 8.1, 7.871645, 7.8, 16.0435, 16.57422, 
    17.12065, 20.44291, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0.9, 7.933333, 10.8, 9.5, 7.9, 7.8, 7.7, 8.15, 8.6, 8.4, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _,
  0.9, 7.933333, 10.8, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _,
  9.5, 9.5, 9.2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _,
  9.1, 7.6, 7.7, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _,
  9.1, 7.6, 7.7, 9.5, 7.9, 7.8, 7.7, 8.15, 8.6, 8.4, 16.57422, 17.12065, 
    20.44291, _, _, _, _, _, _, _, _, _, _, _, _, _,
  9.1, 7.6, 7.7, 9.5, 7.9, 7.8, 7.7, 8.15, 8.6, 8.4, 16.57422, 17.12065, 
    20.44291, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 7.433333, 9.8, 7.1, 8.5, 7.712573, 7, 8.78385, 10.2, 10.3, _, 9.68421, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 7.433333, 9.8, 7.1, 8.5, 7.712573, 7, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 7.433333, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _,
  _, 7.433333, 9.8, 7.1, 8.5, 7.712573, 7, 8.78385, 10.2, 10.3, _, 9.68421, 
    20.44291, _, _, _, _, _, _, _, _, _, _, _, _, _,
  9.5, 7.9, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  9.5, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  1.1, 2.3, 8.7, 8.4, 8.8, 9.260345, 9.6, 9.806979, 9.9, 9.8, _, 9.15, 7.9, 
    _, _, _, _, _, _, _, _, _, _, _, _, _,
  9.5, 9.5, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  9.5, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  9.5, 9.5, 8.7, 8.4, 8.8, 9.260345, 9.6, 9.806979, 9.9, 9.8, _, 9.15, 7.9, 
    _, _, _, _, _, _, _, _, _, _, _, _, _,
  9.5, 9.5, 8.7, 8.4, 8.8, 9.260345, 9.6, 9.806979, 9.9, 9.8, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _,
  9.5, 9.5, 8.7, 8.4, 8.8, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _,
  9.5, 9.5, 8.7, 8.4, 8.8, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _,
  0.1, 0.2, 0.1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _,
  4.8, 2.8, 2.9, 2.2, 3, 1.8, 4.4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _,
  4.8, 2.8, 2.9, 2.2, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _,
  4.8, 2.8, 2.9, 2.2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _,
  7.1, 9.9, 9.433333, 8.966666, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _,
  7.1, 9.9, 9.433333, 8.966666, _, 1.8, 4.4, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _,
  0.6, 2.3, 7.8, 10.4, 8.6, 8.8, 9, 10.24127, 12.1, 9.2, _, 9.25, 9.3, 
    9.8375, 10.7, _, _, _, _, _, _, _, _, _, _, _,
  0.6, 2.3, 7.8, 10.4, 8.6, 8.8, 9, 10.24127, 12.1, 9.2, _, 9.25, 9.3, _, _, 
    _, _, _, _, _, _, _, _, _, _, _,
  0.6, 2.3, 7.8, 10.4, 8.6, 8.8, 9, 10.24127, 12.1, 9.2, _, 9.25, 9.3, 
    9.8375, 10.7, _, _, _, _, _, _, _, _, _, _, _,
  0.6, 2.3, 7.8, 10.4, 8.6, 8.8, 9, 10.24127, 12.1, 9.2, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _,
  0.6, 2.3, 7.8, 10.4, 8.6, 8.8, 9, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _,
  0.6, 2.3, 7.8, 10.4, 8.6, 8.8, 9, 10.24127, 12.1, 9.2, _, 9.25, 9.3, 
    9.8375, _, _, _, _, _, _, _, _, _, _, _, _,
  0.6, 2.3, 7.8, 10.4, 8.6, 8.8, 9, 10.24127, 12.1, 9.2, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _,
  4.2, 6, 4.7, 4, 4.1, 3.1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _,
  4.2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  4.2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  4.2, 6, 4.7, 4, 4.1, 3.1, _, 10.24127, 12.1, 9.2, _, 9.25, 9.3, 9.8375, 
    10.7, _, _, _, _, _, _, _, _, _, _, _,
  4.2, 6, 4.7, 4, 4.1, 3.1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _,
  4.2, 6, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  4.2, 6, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  4.2, 6, 4.7, 4, 4.1, 3.1, _, 10.24127, 12.1, 9.2, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _,
  2.3, 5.3, 9.9, 7.9, 9.1, 9, 8.9, 8.318415, 7.6, 8, _, 8.924999, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _,
  2.3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  2.3, 5.3, 9.9, 7.9, 9.1, 9, 8.9, 8.318415, 7.6, 8, _, 8.924999, 9.3, 
    9.8375, 10.7, _, _, _, _, _, _, _, _, _, _, _,
  2.3, 5.3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  2.3, 5.3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  2.3, 5.3, 9.9, 7.9, 9.1, 9, 8.9, 8.318415, 7.6, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _,
  2.3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  2.3, 5.3, 9.9, 7.9, 9.1, 9, 8.9, 8.318415, 7.6, 8, _, 8.924999, 9.3, 
    9.8375, 10.7, _, _, _, _, _, _, _, _, _, _, _,
  _, 0.09000001, 0.1, 0.1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 0.09000001, 0.1, 0.1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _,
  _, 0.09000001, 0.1, 0.1, 9.1, 9, 8.9, 8.318415, 7.6, 8, _, 8.924999, 9.3, 
    9.8375, 10.7, _, _, _, _, _, _, _, _, _, _, _,
  _, 0.09000001, 0.1, 0.1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _,
  _, 0.09000001, 0.1, 0.1, 9.1, 9, 8.9, 8.318415, 7.6, 8, _, 8.924999, 9.3, 
    9.8375, 10.7, _, _, _, _, _, _, _, _, _, _, _,
  3.8, 4.3, 7.5, 6, 7.5, 7.4, 7.3, 6.834855, 6.2, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _,
  3.8, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  3.8, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  3.8, 4.3, 7.5, 6, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _,
  0.2, 0.1103896, 0.1, 0.1, 0.48, 1.7, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _,
  0.2, 0.1103896, 0.1, 0.1, 0.48, 1.7, 7.3, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _,
  5.9, 8.8, 6.6, 7.9, 6.8, 7.251298, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _,
  5.9, 8.8, 6.6, 7.9, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _,
  5.9, 8.8, 6.6, 7.9, 6.8, 7.251298, 7.3, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _,
  5.9, 8.8, 6.6, 7.9, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _,
  5.9, 8.8, 6.6, 7.9, 6.8, 7.251298, 7.3, 6.834855, 6.2, 8, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _,
  5.9, 8.8, 6.6, 7.9, 6.8, 7.251298, 7.3, 6.834855, 6.2, 8, _, 8.924999, 9.3, 
    9.8375, 10.7, _, _, _, _, _, _, _, _, _, _, _,
  5.9, 8.8, 6.6, 7.9, 6.8, 7.251298, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _,
  5.9, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  5.9, 8.8, 6.6, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _,
  5.9, 8.8, 6.6, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _,
  2.9, 4.6, 5.6, 5.8, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _,
  2.9, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  2.9, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  2.9, 4.6, 5.6, 5.8, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _,
  2.9, 4.6, 5.6, 5.8, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _,
  2.9, 4.6, 5.6, 5.8, 6.8, 7.251298, 7.3, 6.834855, 6.2, 8, _, 8.924999, 9.3, 
    9.8375, 10.7, _, _, _, _, _, _, _, _, _, _, _,
  0.2, 0.02933333, _, _, 0.8535355, 3.445597, _, 11.52235, _, 13.7, 14.24026, 
    14.46415, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  13.8, 11.8, 11.7, 7.2, 5.9, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _,
  13.8, 11.8, 11.7, 7.2, 5.9, 3.445597, _, 11.52235, _, 13.7, 14.24026, 
    14.46415, 9.3, 9.8375, 10.7, _, _, _, _, _, _, _, _, _, _, _,
  13.8, 11.8, 11.7, 7.2, 5.9, 3.445597, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _,
  13.8, 11.8, 11.7, 7.2, 5.9, 3.445597, _, 11.52235, _, 13.7, 14.24026, 
    14.46415, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  13.8, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  13.8, 11.8, 11.7, 7.2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _,
  13.8, 11.8, 11.7, 7.2, 5.9, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _,
  0.2, 0.1158852, 0.04085704, 0.005263157, 0.3, 3.8, 8, 7.871645, 7.8, 
    16.0435, 16.57422, 17.12065, 20.44291, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  0.2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  0.2, 0.1158852, 0.04085704, 0.005263157, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _,
  0.2, 0.1158852, 0.04085704, 0.005263157, 0.3, 3.8, 8, 7.871645, 7.8, 
    16.0435, 16.57422, 17.12065, 20.44291, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  0.2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  0.2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  0.2, 0.1158852, 0.04085704, 0.005263157, 0.3, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _,
  0.2, 0.1158852, 0.04085704, 0.005263157, 0.3, 3.8, 8, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _,
  0.2, 0.1158852, 0.04085704, 0.005263157, 0.3, 3.8, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _,
  0.2, 0.1158852, 0.04085704, 0.005263157, 0.3, 3.8, 8, 7.871645, 7.8, 
    16.0435, 16.57422, 17.12065, 20.44291, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  0.2, 0.1158852, 0.04085704, 0.005263157, 0.3, 3.8, 8, 7.871645, 7.8, 
    16.0435, 16.57422, 17.12065, 20.44291, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  0.2, 0.1158852, 0.04085704, 0.005263157, 0.3, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _,
  0.2, 0.1158852, 0.04085704, 0.005263157, 0.3, 3.8, 8, 7.871645, 7.8, 
    16.0435, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0.2, 0.1158852, 0.04085704, 0.005263157, 0.3, 3.8, 8, 7.871645, 7.8, 
    16.0435, 16.57422, 17.12065, 20.44291, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  7.9, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  14.5, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  14.5, 0.1158852, 0.04085704, 0.005263157, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _,
  11.5, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  11.5, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  7.5, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  7.5, 0.1158852, 0.04085704, 0.005263157, 0.3, 3.8, 8, 7.871645, 7.8, 
    16.0435, 16.57422, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  8.6, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  6.6, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  6.6, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  6.9, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _ ;

 Nitrate_sigfigs =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4, 4, 4, 4, 4, 4, 4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4, 4, 4, 4, 4, 4, 4, 2, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4, 4, 4, 4, 4, 4, 4, 2, 2, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4, 4, 4, 4, 4, 4, 4, 2, 2, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4, 4, 4, 4, 4, 4, 4, 2, 2, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4, 4, 4, 4, 4, 4, 4, 2, 2, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4, 4, 4, 4, 4, 4, 4, 2, 2, 3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, 2, 4, 4, 2, 2, 3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, 2, 4, 4, 2, 2, 3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, 2, 4, 4, 2, 2, 3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, 2, 4, 4, 2, 2, 3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, 2, 4, 4, 2, 2, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, 2, 4, 4, 2, 2, 3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, 2, 4, 4, 2, 2, 3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, 2, 4, 4, 2, 2, 3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, 2, 4, 4, 2, 2, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, 2, 4, 4, 2, 2, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, 2, 4, 4, 2, 2, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, 2, 4, 4, 2, 2, 3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, 2, 4, 4, 2, 2, 3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, 2, 4, 4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, 2, 4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, 2, 2, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, 2, 2, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, 2, 2, 3, 2, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, 2, 2, 3, 2, 2, 2, 2, 2, 3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, 2, 2, 3, 2, 2, 2, 2, 2, 3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, 2, 2, 3, 2, 2, 2, 2, 2, 3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, 2, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, 2, 2, 3, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, 2, 2, 3, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, 2, 2, 3, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, 2, 2, 3, 2, 2, 2, 2, 2, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, 2, 2, 3, 2, 2, 2, 2, 2, 3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, 2, 3, 2, 2, 2, 2, 2, 2, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, 2, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 1, 2, 2, 2, 2, 2, 2, 3, 3, _, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 1, 2, 2, 2, 2, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 1, 2, 2, 2, 2, 2, 2, 3, 3, _, 2, 3, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, 2, 2, 2, 2, 2, 2, _, 2, 2, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, 2, 2, 2, 2, 2, 2, _, 2, 2, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, 2, 2, 2, 2, 2, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, 1, 1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, 2, 2, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, _, 2, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, 2, 2, 3, 2, 2, 2, 3, 3, 2, _, 2, 2, 2, 3, _, _, _, _, _, _, _, _, _, _, _,
  1, 2, 2, 3, 2, 2, 2, 3, 3, 2, _, 2, 2, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, 2, 2, 3, 2, 2, 2, 3, 3, 2, _, 2, 2, 2, 3, _, _, _, _, _, _, _, _, _, _, _,
  1, 2, 2, 3, 2, 2, 2, 3, 3, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, 2, 2, 3, 2, 2, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, 2, 2, 3, 2, 2, 2, 3, 3, 2, _, 2, 2, 2, _, _, _, _, _, _, _, _, _, _, _, _,
  1, 2, 2, 3, 2, 2, 2, 3, 3, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, 2, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, 2, 2, _, 3, 3, 2, _, 2, 2, 2, 3, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, 2, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, 2, 2, _, 3, 3, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, 2, 2, 2, 2, 2, 2, _, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, 2, 2, 2, 2, 2, 2, _, 2, 2, 2, 3, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, 2, 2, 2, 2, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, 2, 2, 2, 2, 2, 2, _, 2, 2, 2, 3, _, _, _, _, _, _, _, _, _, _, _,
  _, 1, 1, 1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 1, 1, 1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 1, 1, 1, 2, 2, 2, 2, 2, 2, _, 2, 2, 2, 3, _, _, _, _, _, _, _, _, _, _, _,
  _, 1, 1, 1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 1, 1, 1, 2, 2, 2, 2, 2, 2, _, 2, 2, 2, 3, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, 2, 2, 2, 2, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, 1, 1, 1, 1, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, 1, 1, 1, 1, 2, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, 2, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, 2, 2, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, 2, 2, 2, 2, 2, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, 2, 2, 2, 2, 2, 2, _, 2, 2, 2, 3, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, 2, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, 2, 2, 2, 2, 2, 2, _, 2, 2, 2, 3, _, _, _, _, _, _, _, _, _, _, _,
  1, 1, _, _, 1, 2, _, 3, _, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, 3, 2, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, 3, 2, 2, 2, _, 3, _, 3, 3, 3, 2, 2, 3, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, 3, 2, 2, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, 3, 2, 2, 2, _, 3, _, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, 3, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, 3, 2, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, 1, 1, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, 1, 1, 1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, 1, 1, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, 1, 1, 1, 1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, 1, 1, 1, 1, 2, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, 1, 1, 1, 1, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, 1, 1, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, 1, 1, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, 1, 1, 1, 1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, 1, 1, 1, 1, 2, 2, 2, 2, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, 1, 1, 1, 1, 2, 2, 2, 2, 3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 1, 1, 1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 1, 1, 1, 1, 2, 2, 2, 2, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 Nitrate_WODflag =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, _, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, _, 0, 0, 0, _, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, _, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _,
  _, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _,
  _, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, _, _, 0, 0, _, 0, _, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, _, 0, _, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, _, 0, _, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 Nitrate_WODprofileflag = _, _, _, _, _, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0 ;

 Nitrate_Original_units =
  "\"ug/l\"    Alternate Nutrient Conversion (use instead of #36)",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "" ;

 pH =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  8.16, 8.12, 8.124302, 8.130274, 8.14, 8.14, 8.14, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _,
  8.16, 8.12, 8.124302, 8.130274, 8.14, 8.14, 8.14, 8.285146, 8.255857, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  8.16, 8.12, 8.124302, 8.130274, 8.14, 8.14, 8.14, 8.285146, 8.255857, 
    8.132226, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  8.16, 8.12, 8.124302, 8.130274, 8.14, 8.14, 8.14, 8.285146, 8.255857, 
    8.132226, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  8.16, 8.12, 8.124302, 8.130274, 8.14, 8.14, 8.14, 8.285146, 8.255857, 
    8.132226, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  8.16, 8.12, 8.124302, 8.130274, 8.14, 8.14, 8.14, 8.285146, 8.255857, 
    8.132226, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  8.16, 8.12, 8.124302, 8.130274, 8.14, 8.14, 8.14, 8.285146, 8.255857, 
    8.132226, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  8.16, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  8.16, 8.12, 8.124302, 8.130274, 8.14, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _,
  8.16, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  8.16, 8.12, 8.124302, 8.130274, 8.14, 8.14, 8.14, 8.285146, 8.255857, 
    8.132226, _, _, _, _, 7.874413, _, _, _, _, _, _, _, _, _, _, _,
  8.16, 8.12, 8.124302, 8.130274, 8.14, 8.14, 8.14, 8.285146, 8.255857, 
    8.132226, _, _, _, _, 7.874413, _, _, _, _, _, _, _, _, _, _, _,
  8.16, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  8.16, 8.12, 8.124302, 8.130274, 8.14, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _,
  8.2, 8.26, 8.253938, 8.25, 8.26, 8.23, 8.2, 8.190795, 8.18, 8.15, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _,
  8.2, 8.26, 8.253938, 8.25, 8.26, 8.23, 8.2, 8.190795, 8.18, 8.15, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _,
  8.2, 8.26, 8.253938, 8.25, 8.26, 8.23, 8.2, 8.190795, 8.18, 8.15, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _,
  8.2, 8.26, 8.253938, 8.25, 8.26, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _,
  8.2, 8.26, 8.253938, 8.25, 8.26, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _,
  8.35, 8.35, 8.35, 8.35, 8.35, 8.35, 8.35, 8.349569, 8.345069, 8.319557, _, 
    _, _, 8.23, _, _, _, _, 8.004101, 7.987364, _, _, _, _, _, _,
  8.35, 8.35, 8.35, 8.35, 8.35, 8.35, 8.35, 8.349569, 8.345069, 8.319557, _, 
    _, _, 8.23, _, _, _, _, _, _, _, _, _, _, _, _,
  8.35, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  8.35, 8.35, 8.35, 8.35, 8.35, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _,
  8.35, 8.35, 8.35, 8.35, 8.35, 8.35, 8.35, 8.349569, 8.345069, 8.319557, _, 
    _, _, 8.23, _, _, _, _, 8.004101, 7.987364, _, _, _, _, _, _,
  8.35, 8.35, 8.35, 8.35, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _,
  8.35, 8.35, 8.35, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _,
  8.35, 8.35, 8.35, 8.35, 8.35, 8.35, 8.35, 8.349569, 8.345069, 8.319557, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  8.35, 8.35, 8.35, 8.35, 8.35, 8.35, 8.35, 8.349569, 8.345069, 8.319557, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  8.35, 8.35, 8.35, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _,
  8.35, 8.35, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _,
  8.35, 8.35, 8.35, 8.35, 8.35, 8.35, 8.35, 8.349569, 8.345069, 8.319557, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  8.35, 8.35, 8.35, 8.35, 8.35, 8.35, 8.35, 8.349569, 8.345069, 8.319557, _, 
    _, _, 8.23, _, _, _, _, 8.004101, 7.987364, _, _, _, _, _, _,
  8.35, 8.35, 8.35, 8.35, 8.35, 8.35, 8.35, 8.349569, 8.345069, 8.319557, _, 
    _, _, 8.23, _, _, _, _, 8.004101, 7.987364, _, _, _, _, _, _,
  8.35, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  8.35, 8.35, 8.35, 8.35, 8.35, 8.35, 8.35, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _,
  8.35, 8.35, 8.35, 8.35, 8.35, 8.35, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _,
  8.35, 8.35, 8.35, 8.35, 8.35, 8.35, 8.35, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _,
  8.35, 8.35, 8.35, 8.35, 8.35, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _,
  8.35, 8.35, 8.35, 8.35, 8.35, 8.35, 8.35, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _,
  8.35, 8.35, 8.35, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _,
  8.35, 8.35, 8.35, 8.35, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _,
  8.35, 8.35, 8.35, 8.35, 8.35, 8.35, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _,
  8.35, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  8.25, 8.248165, 8.244131, 8.237785, 8.218978, 8.19, 8.103258, _, 8.079584, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  8.25, 8.248165, 8.244131, 8.237785, 8.218978, 8.19, 8.103258, _, 8.079584, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  8.25, 8.248165, 8.244131, 8.237785, 8.218978, 8.19, 8.103258, _, 8.079584, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  8.25, 8.248165, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _,
  8.25, 8.248165, 8.244131, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _,
  8.25, 8.248165, 8.244131, 8.237785, 8.218978, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _,
  8.25, 8.248165, 8.244131, 8.237785, 8.218978, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _,
  8.25, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  8.25, 8.248165, 8.244131, 8.237785, 8.218978, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _,
  8.25, 8.248165, 8.244131, 8.237785, 8.218978, 8.19, 8.103258, _, 8.079584, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  8.25, 8.248165, 8.244131, 8.237785, 8.218978, 8.19, 8.103258, _, 8.079584, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  8.25, 8.248165, 8.244131, 8.237785, 8.218978, 8.19, 8.103258, _, 8.079584, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  8.25, 8.248165, 8.244131, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _,
  8.25, 8.248165, 8.244131, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _,
  8.25, 8.248165, 8.244131, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _,
  8.38, 8.368642, 8.35843, 8.349365, 8.334339, 8.322472, 8.320991, 8.328163, 
    8.324529, 8.31, _, _, _, _, _, _, _, _, 8.025373, _, _, _, _, _, _, _,
  8.38, 8.368642, 8.35843, 8.349365, 8.334339, 8.322472, 8.320991, 8.328163, 
    8.324529, 8.31, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  8.38, 8.368642, 8.35843, 8.349365, 8.334339, 8.322472, 8.320991, 8.328163, 
    8.324529, 8.31, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  8.38, 8.368642, 8.35843, 8.349365, 8.334339, 8.322472, 8.320991, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  8.38, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  8.38, 8.368642, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _,
  8.38, 8.368642, 8.35843, 8.349365, 8.334339, 8.322472, 8.320991, 8.328163, 
    8.324529, 8.31, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  8.38, 8.368642, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _,
  8.38, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  8.38, 8.368642, 8.35843, 8.349365, 8.334339, 8.322472, 8.320991, 8.328163, 
    8.324529, 8.31, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  8.38, 8.368642, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _,
  8.38, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  8.38, 8.368642, 8.35843, 8.349365, 8.334339, 8.322472, 8.320991, 8.328163, 
    8.324529, 8.31, _, _, _, _, _, _, _, _, 8.025373, _, _, _, _, _, _, _,
  8.38, 8.368642, 8.35843, 8.349365, 8.334339, 8.322472, 8.320991, 8.328163, 
    8.324529, 8.31, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  8.38, 8.368642, 8.35843, 8.349365, 8.334339, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _,
  8.38, 8.368642, 8.35843, 8.349365, 8.334339, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _,
  8.38, 8.368642, 8.35843, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _,
  8.38, 8.368642, 8.35843, 8.349365, 8.334339, 8.322472, 8.320991, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  8.38, 8.368642, 8.35843, 8.349365, 8.334339, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _,
  8.38, 8.368642, 8.35843, 8.349365, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _,
  8.38, 8.368642, 8.35843, 8.349365, 8.334339, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _,
  8.38, 8.368642, 8.35843, 8.349365, 8.334339, 8.322472, 8.320991, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  8.38, 8.368642, 8.35843, 8.349365, 8.334339, 8.322472, 8.320991, 8.328163, 
    8.324529, 8.31, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  8.38, 8.368642, 8.35843, 8.349365, 8.334339, 8.322472, 8.320991, 8.328163, 
    8.324529, 8.31, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  8.38, 8.368642, 8.35843, 8.349365, 8.334339, 8.322472, 8.320991, 8.328163, 
    8.324529, 8.31, _, _, _, _, _, _, _, _, 8.025373, _, _, _, _, _, _, _,
  8.38, 8.368642, 8.35843, 8.349365, 8.334339, 8.322472, 8.320991, 8.328163, 
    8.324529, 8.31, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  8.38, 8.368642, 8.35843, 8.349365, 8.334339, 8.322472, 8.320991, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  8.38, 8.368642, 8.35843, 8.349365, 8.334339, 8.322472, 8.320991, 8.328163, 
    8.324529, 8.31, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  8.38, 8.368642, 8.35843, 8.349365, 8.334339, 8.322472, 8.320991, 8.328163, 
    8.324529, 8.31, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  8.38, 8.368642, 8.35843, 8.349365, 8.334339, 8.322472, 8.320991, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  8.38, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  8.38, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  8.33, 8.33, 8.33, 8.33, 8.329787, 8.325279, 8.320051, 8.326613, 8.329792, 
    8.318052, _, _, _, _, _, _, _, 8.093211, _, _, _, _, _, _, _, _,
  8.33, 8.33, 8.33, 8.33, 8.329787, 8.325279, 8.320051, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _,
  8.33, 8.33, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _,
  8.33, 8.33, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _,
  8.33, 8.33, 8.33, 8.33, 8.329787, 8.325279, 8.320051, 8.326613, 8.329792, 
    8.318052, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  8.33, 8.33, 8.33, 8.33, 8.329787, 8.325279, 8.320051, 8.326613, 8.329792, 
    8.318052, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  8.33, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  8.33, 8.33, 8.33, 8.33, 8.329787, 8.325279, 8.320051, 8.326613, 8.329792, 
    8.318052, _, _, _, _, _, _, _, 8.093211, _, _, _, _, _, _, _, _,
  8.33, 8.33, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _,
  8.33, 8.33, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _,
  8.33, 8.33, 8.33, 8.33, 8.329787, 8.325279, 8.320051, 8.326613, 8.329792, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  8.33, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  8.33, 8.33, 8.33, 8.33, 8.329787, 8.325279, 8.320051, 8.326613, 8.329792, 
    8.318052, _, _, _, _, _, _, _, 8.093211, _, _, _, _, _, _, _, _,
  8.33, 8.33, 8.33, 8.33, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _,
  8.33, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  8.33, 8.33, 8.33, 8.33, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _,
  8.26, 8.31, 8.30084, 8.292715, 8.29, 8.27, 8.26, 8.2535, 8.25, 8.25, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  8.26, 8.31, 8.30084, 8.292715, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _,
  8.26, 8.31, 8.30084, 8.292715, 8.29, 8.27, 8.26, 8.2535, 8.25, 8.25, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  8.26, 8.31, 8.30084, 8.292715, 8.29, 8.27, 8.26, 8.2535, 8.25, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _,
  8.26, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  8.26, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  8.26, 8.31, 8.30084, 8.292715, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _,
  8.26, 8.31, 8.30084, 8.292715, 8.29, 8.27, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _,
  8.26, 8.31, 8.30084, 8.292715, 8.29, 8.27, 8.26, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _,
  8.26, 8.31, 8.30084, 8.292715, 8.29, 8.27, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _,
  8.26, 8.31, 8.30084, 8.292715, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _,
  8.26, 8.31, 8.30084, 8.292715, 8.29, 8.27, 8.26, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _,
  8.26, 8.31, 8.30084, 8.292715, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _,
  8.26, 8.31, 8.30084, 8.292715, 8.29, 8.27, 8.26, 8.2535, 8.25, 8.25, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  8.25, 8.253802, 8.25759, 8.261366, 8.268879, 8.278169, 8.287357, 8.299107, 
    8.314335, 8.32, 8.310881, _, _, _, _, _, _, _, 8.010458, 7.982935, _, _, 
    _, _, _, _,
  8.25, 8.253802, 8.25759, 8.261366, 8.268879, 8.278169, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _,
  8.25, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  8.25, 8.253802, 8.25759, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _,
  8.25, 8.253802, 8.25759, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _,
  8.25, 8.253802, 8.25759, 8.261366, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _,
  8.25, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  8.25, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  8.25, 8.253802, 8.25759, 8.261366, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _,
  8.25, 8.253802, 8.25759, 8.261366, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _,
  8.25, 8.253802, 8.25759, 8.261366, 8.268879, 8.278169, 8.287357, 8.299107, 
    8.314335, 8.32, 8.310881, _, _, _, _, _, _, _, 8.010458, 7.982935, _, _, 
    _, _, _, _,
  8.25, 8.253802, 8.25759, 8.261366, 8.268879, 8.278169, 8.287357, 8.299107, 
    8.314335, 8.32, 8.310881, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  8.25, 8.253802, 8.25759, 8.261366, 8.268879, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _,
  8.25, 8.253802, 8.25759, 8.261366, 8.268879, 8.278169, 8.287357, 8.299107, 
    8.314335, 8.32, 8.310881, _, _, _, _, _, _, _, 8.010458, 7.982935, _, _, 
    _, _, _, _,
  8.25, 8.253802, 8.25759, 8.261366, 8.268879, 8.278169, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _,
  8.25, 8.253802, 8.25759, 8.261366, 8.268879, 8.278169, 8.287357, 8.299107, 
    8.314335, 8.32, 8.310881, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  8.25, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  8.25, 8.253802, 8.25759, 8.261366, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _,
  8.25, 8.253802, 8.25759, 8.261366, 8.268879, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _,
  8.25, 8.253802, 8.25759, 8.261366, 8.268879, 8.278169, 8.287357, 8.299107, 
    8.314335, 8.32, 8.310881, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  8.25, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  8.25, 8.253802, 8.25759, 8.261366, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _,
  8.27, 8.27811, 8.284187, 8.288229, 8.289017, 8.280513, 8.293255, 8.3, 8.3, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  8.27, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  8.27, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  8.27, 8.27811, 8.284187, 8.288229, 8.289017, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _,
  8.27, 8.27811, 8.284187, 8.288229, 8.289017, 8.280513, 8.293255, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  8.27, 8.27811, 8.284187, 8.288229, 8.289017, 8.280513, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _,
  8.27, 8.28, 8.274824, 8.24, 8.241568, 8.267008, 8.288636, 8.285146, 
    8.255857, 8.132226, _, _, _, _, 7.874413, _, _, _, _, _, _, _, _, _, _, _,
  8.27, 8.28, 8.274824, 8.24, 8.241568, 8.267008, 8.288636, 8.285146, 
    8.255857, 8.132226, _, _, _, _, 7.874413, _, _, _, _, _, _, _, _, _, _, _,
  8.27, 8.28, 8.274824, 8.24, 8.241568, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _,
  8.27, 8.28, 8.274824, 8.24, 8.241568, 8.267008, 8.288636, 8.285146, 
    8.255857, 8.132226, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  8.27, 8.28, 8.274824, 8.24, 8.241568, 8.267008, 8.288636, 8.285146, 
    8.255857, 8.132226, _, _, _, _, 7.874413, _, _, _, _, _, _, _, _, _, _, _,
  8.27, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  8.27, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  8.27, 8.28, 8.274824, 8.24, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _,
  8.27, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  8.27, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  8.27, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  8.27, 8.28, 8.274824, 8.24, 8.241568, 8.267008, 8.288636, 8.285146, 
    8.255857, 8.132226, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  8.27, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  8.27, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  8.27, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  8.27, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _ ;

 pH_sigfigs =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, 3, 3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, 3, 3, 3, 3, 3, 4, 4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, 3, 3, 3, 3, 3, 4, 4, 4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, 3, 3, 3, 3, 3, 4, 4, 4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, 3, 3, 3, 3, 3, 4, 4, 4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, 3, 3, 3, 3, 3, 4, 4, 4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, 3, 3, 3, 3, 3, 4, 4, 4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, 3, 3, 3, 3, 3, 4, 4, 4, _, _, _, _, 4, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, 3, 3, 3, 3, 3, 4, 4, 4, _, _, _, _, 4, _, _, _, _, _, _, _, _, _, _, _,
  3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, 3, 3, 3, 3, 3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, 3, 3, 3, 3, 3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, 3, 3, 3, 3, 3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, 3, 3, 3, 3, 3, 3, 3, 3, 3, _, _, _, 3, _, _, _, _, 3, 3, _, _, _, _, _, _,
  1, 3, 3, 3, 3, 3, 3, 3, 3, 3, _, _, _, 3, _, _, _, _, _, _, _, _, _, _, _, _,
  1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, 3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, 3, 3, 3, 3, 3, 3, 3, 3, 3, _, _, _, 3, _, _, _, _, 3, 3, _, _, _, _, _, _,
  1, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, 3, 3, 3, 3, 3, 3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, 3, 3, 3, 3, 3, 3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, 3, 3, 3, 3, 3, 3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, 3, 3, 3, 3, 3, 3, 3, 3, 3, _, _, _, 3, _, _, _, _, 3, 3, _, _, _, _, _, _,
  1, 3, 3, 3, 3, 3, 3, 3, 3, 3, _, _, _, 3, _, _, _, _, 3, 3, _, _, _, _, _, _,
  1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, 3, 3, 3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, 3, 3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, 3, 3, 3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, 3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, 3, 3, 3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, 3, 3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, 3, 3, 3, 3, 3, 3, _, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, 3, 3, 3, 3, 3, 3, _, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, 3, 3, 3, 3, 3, 3, _, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, 3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, 3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, 3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, 3, 3, 3, 3, 3, 3, _, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, 3, 3, 3, 3, 3, 3, _, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, 3, 3, 3, 3, 3, 3, _, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, 3, 3, 3, 3, 3, 3, 3, 3, 3, _, _, _, _, _, _, _, _, 3, _, _, _, _, _, _, _,
  1, 3, 3, 3, 3, 3, 3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, 3, 3, 3, 3, 3, 3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, 3, 3, 3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, 3, 3, 3, 3, 3, 3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, 3, 3, 3, 3, 3, 3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, 3, 3, 3, 3, 3, 3, 3, 3, 3, _, _, _, _, _, _, _, _, 3, _, _, _, _, _, _, _,
  1, 3, 3, 3, 3, 3, 3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, 3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, 3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, 3, 3, 3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, 3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, 3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, 3, 3, 3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, 3, 3, 3, 3, 3, 3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, 3, 3, 3, 3, 3, 3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, 3, 3, 3, 3, 3, 3, 3, 3, 3, _, _, _, _, _, _, _, _, 3, _, _, _, _, _, _, _,
  1, 3, 3, 3, 3, 3, 3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, 3, 3, 3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, 3, 3, 3, 3, 3, 3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, 3, 3, 3, 3, 3, 3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, 3, 3, 3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, 3, 3, 3, 3, 3, 3, 3, 3, 3, _, _, _, _, _, _, _, 3, _, _, _, _, _, _, _, _,
  1, 3, 3, 3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, 3, 3, 3, 3, 3, 3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, 3, 3, 3, 3, 3, 3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, 3, 3, 3, 3, 3, 3, 3, 3, 3, _, _, _, _, _, _, _, 3, _, _, _, _, _, _, _, _,
  1, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, 3, 3, 3, 3, 3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, 3, 3, 3, 3, 3, 3, 3, 3, 3, _, _, _, _, _, _, _, 3, _, _, _, _, _, _, _, _,
  1, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, 3, 3, 3, 3, 3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, 3, 3, 3, 3, 3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, 3, 3, 3, 3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, 3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, 3, 3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, 3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, 3, 3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, 3, 3, 3, 3, 3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, _, _, _, _, _, _, _, 3, 3, _, _, _, _, _, _,
  1, 3, 3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, _, _, _, _, _, _, _, 3, 3, _, _, _, _, _, _,
  1, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, 3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, _, _, _, _, _, _, _, 3, 3, _, _, _, _, _, _,
  1, 3, 3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, 3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, 3, 3, 3, 3, 3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, 3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, 3, 3, 3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, 3, 3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4, 4, 4, 4, 4, 4, 4, 4, 4, 4, _, _, _, _, 4, _, _, _, _, _, _, _, _, _, _, _,
  4, 4, 4, 4, 4, 4, 4, 4, 4, 4, _, _, _, _, 4, _, _, _, _, _, _, _, _, _, _, _,
  4, 4, 4, 4, 4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4, 4, 4, 4, 4, 4, 4, 4, 4, 4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4, 4, 4, 4, 4, 4, 4, 4, 4, 4, _, _, _, _, 4, _, _, _, _, _, _, _, _, _, _, _,
  4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4, 4, 4, 4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4, 4, 4, 4, 4, 4, 4, 4, 4, 4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 pH_WODflag =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, 0, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, 0, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, 0, _, _, _, _, 0, 0, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, 0, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, 0, _, _, _, _, 0, 0, _, _, _, _, _, _,
  0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, 0, _, _, _, _, 0, 0, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, 0, _, _, _, _, 0, 0, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, 0, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, 0, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, 0, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, 0, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, 0, _, _, _, _, _, _, _, _,
  0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, 0, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, 0, 0, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, 0, 0, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, 0, 0, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, 0, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, 0, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, 0, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 pH_WODprofileflag = _, _, _, _, _, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0 ;

 Ammonia =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1.4, 3.1, 3.7, 2.6, 2.6, 2.728571, 3, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _,
  1.4, 3.1, 3.7, 2.6, 2.6, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _,
  1.4, 3.1, 3.7, 2.6, 2.6, 2.728571, 3, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _,
  1.4, 3.1, 3.7, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _,
  1.4, 3.1, 3.7, 2.6, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _,
  1.4, 1.8, 3.3, 1.8, 0.5, 2.3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _,
  1.4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  1.4, 1.8, 3.3, 1.8, 0.5, 2.3, 3, 0.6003202, _, 0.3, 0.3697152, 0.4, 1.4, 
    1.1875, 0.4, _, _, _, _, _, _, _, _, _, _, _,
  1.4, 1.8, 3.3, 1.8, 0.5, 2.3, 3, 0.6003202, _, 0.3, 0.3697152, 0.4, 1.4, 
    1.1875, 0.4, _, _, _, _, _, _, _, _, _, _, _,
  1.4, 1.8, 3.3, 1.8, 0.5, 2.3, 3, 0.6003202, _, 0.3, 0.3697152, 0.4, 1.4, 
    1.1875, 0.4, _, _, _, _, _, _, _, _, _, _, _,
  1.4, 1.8, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  1.4, 1.8, 3.3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _,
  1.4, 1.8, 3.3, 1.8, 0.5, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _,
  1.4, 1.8, 3.3, 1.8, 0.5, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _,
  1.4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  1.4, 1.8, 3.3, 1.8, 0.5, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _,
  1.4, 1.8, 3.3, 1.8, 0.5, 2.3, 3, 0.6003202, _, 0.3, 0.3697152, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _,
  1.4, 1.8, 3.3, 1.8, 0.5, 2.3, 3, 0.6003202, _, 0.3, 0.3697152, 0.4, 1.4, 
    1.1875, 0.4, _, _, _, _, _, _, _, _, _, _, _,
  0.7, 1.7, 1.1, 0.4, 0.7, 0.7167073, 0.8, 0.9659172, 1.2, 0.8, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _,
  0.7, 1.7, 1.1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _,
  0.7, 1.7, 1.1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _,
  0.7, 1.7, 1.1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _,
  0.7, 1.7, 1.1, 0.4, 0.7, 0.7167073, 0.8, 0.9659172, 1.2, 0.8, 0.3697152, 
    0.4, 1.4, 1.1875, 0.4, _, _, _, _, _, _, _, _, _, _, _,
  0.7, 1.7, 1.1, 0.4, 0.7, 0.7167073, 0.8, 0.9659172, 1.2, 0.8, 0.3697152, 
    0.4, 1.4, 1.1875, 0.4, _, _, _, _, _, _, _, _, _, _, _,
  0.6, 0.5, 0.2, 0.5, 0.5, 0.8147652, 1.2, 1.02561, 0.9, 1.4, _, 1.347368, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _,
  0.6, 0.5, 0.2, 0.5, 0.5, 0.8147652, 1.2, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _,
  0.6, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  0.6, 0.5, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  0.6, 0.5, 0.2, 0.5, 0.5, 0.8147652, 1.2, 1.02561, 0.9, 1.4, _, 1.347368, 
    1.4, 1.1875, 0.4, _, _, _, _, _, _, _, _, _, _, _,
  0.6, 0.5, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  0.6, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  0.8, 0.4, 0.5, 0.3, 1.3, 1.2, 1.1, 0.7266423, 0.2, 0.8, _, 0.85, 0.9, _, _, 
    _, _, _, _, _, _, _, _, _, _, _,
  0.8, 0.4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  0.8, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  0.8, 0.4, 0.5, 0.3, 1.3, 1.2, 1.1, 0.7266423, 0.2, 0.8, _, 0.85, 0.9, 
    1.1875, 0.4, _, _, _, _, _, _, _, _, _, _, _,
  0.8, 0.4, 0.5, 0.3, 1.3, 1.2, 1.1, 0.7266423, 0.2, 0.8, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _,
  0.8, 0.4, 0.5, 0.3, 1.3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _,
  0.8, 0.4, 0.5, 0.3, 1.3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _,
  1.7, 0.6, 0.5272727, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _,
  1.7, 0.6, 0.5272727, 0.3, 1.3, 1.2, 1.1, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _,
  1.7, 0.6, 0.5272727, 0.3, 1.3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _,
  1.7, 0.6, 0.5272727, 0.3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _,
  1.7, 0.6, 0.5272727, 0.3, 1.3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _,
  1.7, 0.6, 0.5272727, 0.3, 1.3, 1.2, 1.1, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _,
  1, 1.3, 1.1, 2, 0.2, 0.2, 0.2, 0.5133145, 1, 0.1, _, 0.75, 1.4, 1.1875, 
    0.4, _, _, _, _, _, _, _, _, _, _, _,
  1, 1.3, 1.1, 2, 0.2, 0.2, 0.2, 0.5133145, 1, 0.1, _, 0.75, 1.4, _, _, _, _, 
    _, _, _, _, _, _, _, _, _,
  1, 1.3, 1.1, 2, 0.2, 0.2, 0.2, 0.5133145, 1, 0.1, _, 0.75, 1.4, 1.1875, 
    0.4, _, _, _, _, _, _, _, _, _, _, _,
  1, 1.3, 1.1, 2, 0.2, 0.2, 0.2, 0.5133145, 1, 0.1, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _,
  1, 1.3, 1.1, 2, 0.2, 0.2, 0.2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _,
  1, 1.3, 1.1, 2, 0.2, 0.2, 0.2, 0.5133145, 1, 0.1, _, 0.75, 1.4, 1.1875, _, 
    _, _, _, _, _, _, _, _, _, _, _,
  1, 1.3, 1.1, 2, 0.2, 0.2, 0.2, 0.5133145, 1, 0.1, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _,
  1, 1.3, 1.1, 2, 0.2, 0.2, 0.2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _,
  1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, 1.3, 1.1, 2, 0.2, 0.2, 0.2, 0.5133145, 1, 0.1, _, 0.75, 1.4, 1.1875, 
    0.4, _, _, _, _, _, _, _, _, _, _, _,
  1, 1.3, 1.1, 2, 0.2, 0.2, 0.2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _,
  1, 1.3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  1, 1.3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  1, 1.3, 1.1, 2, 0.2, 0.2, 0.2, 0.5133145, 1, 0.1, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _,
  0.7, 1.1, 0.2, 0.7, 1.8, 1.440366, 1.1, 0.8459134, 0.7, 0.8, _, 1.072369, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0.7, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  0.7, 1.1, 0.2, 0.7, 1.8, 1.440366, 1.1, 0.8459134, 0.7, 0.8, _, 1.072369, 
    1.4, 1.1875, 0.4, _, _, _, _, _, _, _, _, _, _, _,
  0.7, 1.1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  0.7, 1.1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  0.7, 1.1, 0.2, 0.7, 1.8, 1.440366, 1.1, 0.8459134, 0.7, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _,
  0.7, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  0.7, 1.1, 0.2, 0.7, 1.8, 1.440366, 1.1, 0.8459134, 0.7, 0.8, _, 1.072369, 
    1.4, 1.1875, 0.4, _, _, _, _, _, _, _, _, _, _, _,
  0.8, 0.64, 0.4227059, 0.6, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _,
  0.8, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  0.8, 0.64, 0.4227059, 0.6, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _,
  0.8, 0.64, 0.4227059, 0.6, 1.8, 1.440366, 1.1, 0.8459134, 0.7, 0.8, _, 
    1.072369, 1.4, 1.1875, 0.4, _, _, _, _, _, _, _, _, _, _, _,
  0.8, 0.64, 0.4227059, 0.6, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _,
  0.8, 0.64, 0.4227059, 0.6, 1.8, 1.440366, 1.1, 0.8459134, 0.7, 0.8, _, 
    1.072369, 1.4, 1.1875, 0.4, _, _, _, _, _, _, _, _, _, _, _,
  0.8, 0.9, 1.2, 0.8, 1.6, 0.8504452, 0.4, 0.7718408, 1, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _,
  0.8, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  0.8, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  0.8, 0.9, 1.2, 0.8, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _,
  1.3, 1.146494, 0.8624626, 0.9777778, 1.511516, 1.8, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _,
  1.3, 1.146494, 0.8624626, 0.9777778, 1.511516, 1.8, 0.4, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, 1, 1.1, 1.2, 0.2, 0.4142857, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _,
  1, 1, 1.1, 1.2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  1, 1, 1.1, 1.2, 0.2, 0.4142857, 0.4, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _,
  1, 1, 1.1, 1.2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  1, 1, 1.1, 1.2, 0.2, 0.4142857, 0.4, 0.7718408, 1, 0.8, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _,
  1, 1, 1.1, 1.2, 0.2, 0.4142857, 0.4, 0.7718408, 1, 0.8, _, 1.072369, 1.4, 
    1.1875, 0.4, _, _, _, _, _, _, _, _, _, _, _,
  1, 1, 1.1, 1.2, 0.2, 0.4142857, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _,
  1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, 1, 1.1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  1, 1, 1.1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  0.5, 0.5, 0.5, 1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _,
  0.5, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  0.5, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  0.5, 0.5, 0.5, 1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _,
  0.5, 0.5, 0.5, 1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _,
  0.5, 0.5, 0.5, 1, 0.2, 0.4142857, 0.4, 0.7718408, 1, 0.8, _, 1.072369, 1.4, 
    1.1875, 0.4, _, _, _, _, _, _, _, _, _, _, _,
  1, 0.6586667, 0.6, 0.6, 0.7841707, 0.8958333, _, 0.6003202, _, 0.3, 
    0.3697152, 0.4, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3.6, 3.6, 3.1, 3.2, 0.7, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _,
  3.6, 3.6, 3.1, 3.2, 0.7, 0.8958333, _, 0.6003202, _, 0.3, 0.3697152, 0.4, 
    1.4, 1.1875, 0.4, _, _, _, _, _, _, _, _, _, _, _,
  3.6, 3.6, 3.1, 3.2, 0.7, 0.8958333, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _,
  3.6, 3.6, 3.1, 3.2, 0.7, 0.8958333, _, 0.6003202, _, 0.3, 0.3697152, 0.4, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3.6, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  3.6, 3.6, 3.1, 3.2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _,
  3.6, 3.6, 3.1, 3.2, 0.7, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _,
  3.6, 3.6, 3.1, 3.2, 0.7, 0.8958333, _, 0.6003202, _, 0.3, 0.3697152, 0.4, 
    1.4, 1.1875, 0.4, _, _, _, _, _, _, _, _, _, _, _,
  3.6, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  3.6, 3.6, 3.1, 3.2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _,
  3.6, 3.6, 3.1, 3.2, 0.7, 0.8958333, _, 0.6003202, _, 0.3, 0.3697152, 0.4, 
    1.4, 1.1875, 0.4, _, _, _, _, _, _, _, _, _, _, _,
  3.6, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  3.6, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  3.6, 3.6, 3.1, 3.2, 0.7, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _,
  3.6, 3.6, 3.1, 3.2, 0.7, 0.8958333, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _,
  3.6, 3.6, 3.1, 3.2, 0.7, 0.8958333, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _,
  3.6, 3.6, 3.1, 3.2, 0.7, 0.8958333, _, 0.6003202, _, 0.3, 0.3697152, 0.4, 
    1.4, 1.1875, 0.4, _, _, _, _, _, _, _, _, _, _, _,
  3.6, 3.6, 3.1, 3.2, 0.7, 0.8958333, _, 0.6003202, _, 0.3, 0.3697152, 0.4, 
    1.4, 1.1875, 0.4, _, _, _, _, _, _, _, _, _, _, _,
  3.6, 3.6, 3.1, 3.2, 0.7, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _,
  3.6, 3.6, 3.1, 3.2, 0.7, 0.8958333, _, 0.6003202, _, 0.3, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _,
  3.6, 3.6, 3.1, 3.2, 0.7, 0.8958333, _, 0.6003202, _, 0.3, 0.3697152, 0.4, 
    1.4, 1.1875, 0.4, _, _, _, _, _, _, _, _, _, _, _,
  3.6, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  3.6, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  3.6, 3.6, 3.1, 3.2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _,
  3.6, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  3.6, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  3.6, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  3.6, 3.6, 3.1, 3.2, 0.7, 0.8958333, _, 0.6003202, _, 0.3, 0.3697152, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _,
  3.6, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  3.6, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  3.6, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  3.6, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _ ;

 Ammonia_sigfigs =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, 2, 2, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, 2, 2, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, 1, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, 1, 2, 2, 1, _, 1, 1, 1, 2, 2, 1, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, 1, 2, 2, 1, _, 1, 1, 1, 2, 2, 1, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, 1, 2, 2, 1, _, 1, 1, 1, 2, 2, 1, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, 1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, 1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, 1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, 1, 2, 2, 1, _, 1, 1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, 1, 2, 2, 1, _, 1, 1, 1, 2, 2, 1, _, _, _, _, _, _, _, _, _, _, _,
  1, 2, 2, 1, 1, 1, 1, 2, 2, 1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, 2, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, 2, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, 2, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, 2, 2, 1, 1, 1, 1, 2, 2, 1, 1, 1, 2, 2, 1, _, _, _, _, _, _, _, _, _, _, _,
  1, 2, 2, 1, 1, 1, 1, 2, 2, 1, 1, 1, 2, 2, 1, _, _, _, _, _, _, _, _, _, _, _,
  1, 1, 1, 1, 1, 1, 2, 2, 1, 2, _, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, 1, 1, 1, 1, 1, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, 1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, 1, 1, 1, 1, 1, 2, 2, 1, 2, _, 2, 2, 2, 1, _, _, _, _, _, _, _, _, _, _, _,
  1, 1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, 1, 1, 1, 2, 2, 2, 1, 1, 1, _, 1, 1, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, 1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, 1, 1, 1, 2, 2, 2, 1, 1, 1, _, 1, 1, 2, 1, _, _, _, _, _, _, _, _, _, _, _,
  1, 1, 1, 1, 2, 2, 2, 1, 1, 1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, 1, 1, 1, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, 1, 1, 1, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, 1, 1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, 1, 1, 1, 2, 2, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, 1, 1, 1, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, 1, 1, 1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, 1, 1, 1, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, 1, 1, 1, 2, 2, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, 1, 1, 1, 1, 2, 1, _, 1, 2, 2, 1, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, 1, 1, 1, 1, 2, 1, _, 1, 2, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, 1, 1, 1, 1, 2, 1, _, 1, 2, 2, 1, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, 1, 1, 1, 1, 2, 1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, 1, 1, 1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, 1, 1, 1, 1, 2, 1, _, 1, 2, 2, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, 1, 1, 1, 1, 2, 1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, 1, 1, 1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, 1, 1, 1, 1, 2, 1, _, 1, 2, 2, 1, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, 1, 1, 1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, 1, 1, 1, 1, 2, 1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, 2, 1, 1, 2, 2, 2, 1, 1, 1, _, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, 2, 1, 1, 2, 2, 2, 1, 1, 1, _, 2, 2, 2, 1, _, _, _, _, _, _, _, _, _, _, _,
  1, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, 2, 1, 1, 2, 2, 2, 1, 1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, 2, 1, 1, 2, 2, 2, 1, 1, 1, _, 2, 2, 2, 1, _, _, _, _, _, _, _, _, _, _, _,
  1, 1, 1, 1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, 1, 1, 1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, 1, 1, 1, 2, 2, 2, 1, 1, 1, _, 2, 2, 2, 1, _, _, _, _, _, _, _, _, _, _, _,
  1, 1, 1, 1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, 1, 1, 1, 2, 2, 2, 1, 1, 1, _, 2, 2, 2, 1, _, _, _, _, _, _, _, _, _, _, _,
  1, 1, 2, 1, 2, 1, 1, 1, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, 1, 2, 1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, 2, 1, 2, 2, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, 2, 1, 2, 2, 2, 1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, 1, 1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, 1, 1, 1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, 1, 1, 1, 1, 2, 1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, 1, 1, 1, 1, 2, 1, _, 2, 2, 2, 1, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, 1, 1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, 1, 1, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, 1, 1, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, 1, 1, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, 1, 1, 2, 1, 1, 1, 1, 2, 1, _, 2, 2, 2, 1, _, _, _, _, _, _, _, _, _, _, _,
  1, 1, 1, 1, 1, 1, _, 1, _, 1, 1, 1, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, 1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, 1, 1, _, 1, _, 1, 1, 1, 2, 2, 1, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, 1, 1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, 1, 1, _, 1, _, 1, 1, 1, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, 1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, 1, 1, _, 1, _, 1, 1, 1, 2, 2, 1, _, _, _, _, _, _, _, _, _, _, _,
  2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, 1, 1, _, 1, _, 1, 1, 1, 2, 2, 1, _, _, _, _, _, _, _, _, _, _, _,
  2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, 1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, 1, 1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, 1, 1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, 1, 1, _, 1, _, 1, 1, 1, 2, 2, 1, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, 1, 1, _, 1, _, 1, 1, 1, 2, 2, 1, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, 1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, 1, 1, _, 1, _, 1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, 1, 1, _, 1, _, 1, 1, 1, 2, 2, 1, _, _, _, _, _, _, _, _, _, _, _,
  2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, 1, 1, _, 1, _, 1, 1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 Ammonia_WODflag =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, _, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, _, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, _, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, _, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, _, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, _, 0, _, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, _, 0, _, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, _, 0, _, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, _, 0, _, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, _, 0, _, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, _, 0, _, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, _, 0, _, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, _, 0, _, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, _, 0, _, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, _, 0, _, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 Chlorophyll =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0.425, 0.604, 0.439, 0.606, 0.444, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _,
  0.425, 0.604, 0.439, 0.606, 0.444, 0.4, 0.1, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _,
  0.425, 0.604, 0.439, 0.606, 0.444, 0.4, 0.1, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _,
  0.425, 0.604, 0.439, 0.606, 0.444, 0.4, 0.1, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _,
  0.425, 0.604, 0.439, 0.606, 0.444, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _,
  0.425, 0.604, 0.439, 0.606, 0.444, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _,
  0.425, 0.604, 0.439, 0.606, 0.444, 0.4, 0.1, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _,
  0.425, 0.604, 0.439, 0.606, 0.444, 0.4, 0.1, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _,
  0.425, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  0.425, 0.604, 0.439, 0.606, 0.444, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _,
  0.425, 0.604, 0.439, 0.606, 0.444, 0.4, 0.1, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _,
  0.425, 0.604, 0.439, 0.606, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _,
  1.1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  1.1, _, _, 0.606, 0.444, 0.4, 0.1, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _,
  1.1, _, _, 0.606, 0.444, 0.4, 0.1, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _,
  1.121, 1.027, 1.316333, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _,
  1.121, 1.027, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _,
  1.121, 1.027, 1.316333, 0.606, 0.444, 0.4, 0.1, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _,
  1.121, 1.027, 1.316333, 0.606, 0.444, 0.4, 0.1, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _,
  1.121, 1.027, 1.316333, 0.606, 0.444, 0.4, 0.1, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _,
  1.121, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  1.121, 1.027, 1.316333, 0.606, 0.444, 0.4, 0.1, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _,
  1.121, 1.027, 1.316333, 0.606, 0.444, 0.4, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _,
  22.3, 21.8, 12.2, 0.4, 0.1, 0.1, 0.1, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _,
  22.3, 21.8, 12.2, 0.4, 0.1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _,
  22.3, 21.8, 12.2, 0.4, 0.1, 0.1, 0.1, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _,
  22.3, 21.8, 12.2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _,
  22.3, 21.8, 12.2, 0.4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _,
  30.2, 17.4, 12.5, 0.6, 0.2, 0.1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _,
  30.2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  30.2, 17.4, 12.5, 0.6, 0.2, 0.1, 0.1, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _,
  30.2, 17.4, 12.5, 0.6, 0.2, 0.1, 0.1, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _,
  30.2, 17.4, 12.5, 0.6, 0.2, 0.1, 0.1, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _,
  30.2, 17.4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _,
  1.7, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  1.7, _, _, 0.6, 0.2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _,
  1.7, _, _, 0.6, 0.2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _,
  1.7, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  0.636, 0.729, 0.431, 0.856, 0.809, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _,
  0.636, 0.729, 0.431, 0.856, 0.809, 0.1, 0.1, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _,
  0.636, 0.729, 0.431, 0.856, 0.809, 0.1, 0.1, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _,
  0.636, 0.729, 0.431, 0.856, 0.809, 0.1, 0.1, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _,
  1.665, 1.582, 1.594, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _,
  1.665, 1.582, 1.594, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _,
  1.665, 1.582, 1.594, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _,
  1.665, 1.582, 1.594, 0.856, 0.809, 0.1, 0.1, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _,
  1.665, 1.582, 1.594, 0.856, 0.809, 0.1, 0.1, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _,
  33.5, 1.8, 0.5, 0.2, 0.2, 0.2, 0.1, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _,
  33.5, 1.8, 0.5, 0.2, 0.2, 0.2, 0.1, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _,
  33.5, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  33.5, 1.8, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _,
  33.5, 1.8, 0.5, 0.2, 0.2, 0.2, 0.1, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _,
  33.5, 1.8, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _,
  33.5, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  33.5, 1.8, 0.5, 0.2, 0.2, 0.2, 0.1, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _,
  33.5, 1.8, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _,
  33.5, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  33.5, 1.8, 0.5, 0.2, 0.2, 0.2, 0.1, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _,
  33.5, 1.8, 0.5, 0.2, 0.2, 0.2, 0.1, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _,
  3.2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  3.2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  3.2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  3.2, _, _, _, _, 0.2, 0.1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _,
  2.759, 2.579, 2.357879, 3.49, 5.042, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _,
  3.203, 3.312, 1.535, 3.025, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _,
  3.203, 3.312, 1.535, 3.025, 5.042, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _,
  3.203, 3.312, 1.535, 3.025, 5.042, 0.2, 0.1, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _,
  24.7, 19, 0.4, 0.3, 0.2, 0.1, 0.1, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _,
  24.7, 19, 0.4, 0.3, 0.2, 0.1, 0.1, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _,
  24.7, 19, 0.4, 0.3, 0.2, 0.1, 0.1, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _,
  24.7, 19, 0.4, 0.3, 0.2, 0.1, 0.1, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _,
  24.7, 19, 0.4, 0.3, 0.2, 0.1, 0.1, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _,
  24.7, 19, 0.4, 0.3, 0.2, 0.1, 0.1, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _,
  24.7, 19, 0.4, 0.3, 0.2, 0.1, 0.1, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _,
  24.7, 19, 0.4, 0.3, 0.2, 0.1, 0.1, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _,
  24.7, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  24.7, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  24.7, 19, 0.4, 0.3, 0.2, 0.1, 0.1, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _,
  24.7, 19, 0.4, 0.3, 0.2, 0.1, 0.1, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _,
  24.7, 19, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  24.7, 19, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  24.7, 19, 0.4, 0.3, 0.2, 0.1, 0.1, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _,
  17.3, 12.3, 0.3, 0.2, 0.2, 0.2, 0.1, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _,
  17.3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  17.3, 12.3, 0.3, 0.2, 0.2, 0.2, 0.1, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _,
  17.3, 12.3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _,
  17.3, 12.3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _,
  17.3, 12.3, 0.3, 0.2, 0.2, 0.2, 0.1, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _,
  17.3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  17.3, 12.3, 0.3, 0.2, 0.2, 0.2, 0.1, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _,
  17.3, 12.3, 0.3, 0.2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _,
  17.3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  2.177, 2.285, 2.085, 1.881, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _,
  2.177, 2.285, 2.085, 1.881, 0.2, 0.2, 0.1, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _,
  0.6, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  0.6, _, _, _, 0.2, 0.2, 0.1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _,
  0.6, _, _, _, 0.2, 0.2, 0.1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _,
  0.6, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  0.6, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  0.597, 0.4083333, 0.2877479, 0.981, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _,
  0.597, 0.4083333, 0.2877479, 0.981, 0.2, 0.2, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _,
  0.597, 0.4083333, 0.2877479, 0.981, 0.2, 0.2, 0.1, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _,
  9.3, 6.7, 3.7, 0.4, 0.3, 0.4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _,
  9.3, 6.7, 3.7, 0.4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _,
  9.3, 6.7, 3.7, 0.4, 0.3, 0.4, 0.1, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _,
  9.3, 6.7, 3.7, 0.4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _,
  9.3, 6.7, 3.7, 0.4, 0.3, 0.4, 0.1, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _,
  9.3, 6.7, 3.7, 0.4, 0.3, 0.4, 0.1, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _,
  9.3, 6.7, 3.7, 0.4, 0.3, 0.4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _,
  9.3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  0.657, 0.575, 1.059, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _,
  0.657, 0.575, 1.059, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _,
  0.657, 0.575, 1.059, 0.4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _,
  0.657, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  0.657, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  0.657, 0.575, 1.059, 0.4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _,
  0.657, 0.575, 1.059, 0.4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _,
  0.657, 0.575, 1.059, 0.4, 0.3, 0.4, 0.1, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _,
  0.657, 0.575, 1.059, 0.4, 0.3, 0.4, 0.1, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _,
  1.4, 1.1, 1, 1.1, 0.3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _,
  1.4, 1.1, 1, 1.1, 0.3, 0.4, 0.1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _,
  1.4, 1.1, 1, 1.1, 0.3, 0.4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _,
  1.4, 1.1, 1, 1.1, 0.3, 0.4, 0.1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _,
  1.4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  1.4, 1.1, 1, 1.1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _,
  1.4, 1.1, 1, 1.1, 0.3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _,
  1.4, 1.1, 1, 1.1, 0.3, 0.4, 0.1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _,
  1.4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  0.28, 0.283, 0.385, 0.99, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _,
  0.28, 0.283, 0.385, 0.99, 0.3, 0.4, 0.1, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _,
  0.28, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  0.28, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  0.59, 0.701, 0.716, 1.67, 2.024, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _,
  0.59, 0.701, 0.716, 1.67, 2.024, 0.4, 0.1, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _,
  0.59, 0.701, 0.716, 1.67, 2.024, 0.4, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _,
  0.59, 0.701, 0.716, 1.67, 2.024, 0.4, 0.1, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _,
  0.59, 0.701, 0.716, 1.67, 2.024, 0.4, 0.1, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _,
  0.59, 0.701, 0.716, 1.67, 2.024, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _,
  0.59, 0.701, 0.716, 1.67, 2.024, 0.4, 0.1, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _,
  0.59, 0.701, 0.716, 1.67, 2.024, 0.4, 0.1, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _,
  0.59, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  0.59, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  0.59, 0.701, 0.716, 1.67, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _,
  0.59, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  3.02, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  3.02, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  3.02, 0.701, 0.716, 1.67, 2.024, 0.4, 0.1, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _,
  3.02, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  3.02, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  3.02, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  3.02, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _ ;

 Chlorophyll_sigfigs =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, 3, 3, 3, 1, 1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, 3, 3, 3, 1, 1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, 3, 3, 3, 1, 1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, 3, 3, 3, 1, 1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, 3, 3, 3, 1, 1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, 3, 3, 3, 1, 1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, _, _, 3, 3, 1, 1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, _, _, 3, 3, 1, 1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4, 4, 4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4, 4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4, 4, 4, 3, 3, 1, 1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4, 4, 4, 3, 3, 1, 1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4, 4, 4, 3, 3, 1, 1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4, 4, 4, 3, 3, 1, 1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4, 4, 4, 3, 3, 1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, 3, 1, 1, 1, 1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, 3, 1, 1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, 3, 1, 1, 1, 1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, 3, 1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, 3, 1, 1, 1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, 3, 1, 1, 1, 1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, 3, 1, 1, 1, 1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, 3, 1, 1, 1, 1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, _, _, 1, 1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, _, _, 1, 1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, 3, 3, 3, 1, 1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, 3, 3, 3, 1, 1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, 3, 3, 3, 1, 1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4, 4, 4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4, 4, 4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4, 4, 4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4, 4, 4, 3, 3, 1, 1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4, 4, 4, 3, 3, 1, 1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 2, 1, 1, 1, 1, 1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 2, 1, 1, 1, 1, 1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 2, 1, 1, 1, 1, 1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 2, 1, 1, 1, 1, 1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 2, 1, 1, 1, 1, 1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 2, 1, 1, 1, 1, 1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, _, _, _, _, 1, 1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4, 4, 4, 4, 4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4, 4, 4, 4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4, 4, 4, 4, 4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4, 4, 4, 4, 4, 1, 1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, 1, 1, 1, 1, 1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, 1, 1, 1, 1, 1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, 1, 1, 1, 1, 1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, 1, 1, 1, 1, 1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, 1, 1, 1, 1, 1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, 1, 1, 1, 1, 1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, 1, 1, 1, 1, 1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, 1, 1, 1, 1, 1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, 1, 1, 1, 1, 1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, 1, 1, 1, 1, 1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, 1, 1, 1, 1, 1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, 1, 1, 1, 1, 1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, 1, 1, 1, 1, 1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, 1, 1, 1, 1, 1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, 1, 1, 1, 1, 1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, 1, 1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4, 4, 4, 4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4, 4, 4, 4, 1, 1, 1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, _, _, _, 1, 1, 1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, _, _, _, 1, 1, 1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, 3, 3, 1, 1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, 3, 3, 1, 1, 1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 1, 1, 1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 1, 1, 1, 1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 1, 1, 1, 1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 1, 1, 1, 1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 1, 1, 1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, 4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, 4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, 4, 1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, 4, 1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, 4, 1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, 4, 1, 1, 1, 1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, 4, 1, 1, 1, 1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, 1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, 1, 1, 1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, 1, 1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, 1, 1, 1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, 1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, 2, 2, 2, 1, 1, 1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, 3, 3, 1, 1, 1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, 3, 4, 4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, 3, 4, 4, 1, 1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, 3, 4, 4, 1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, 3, 4, 4, 1, 1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, 3, 4, 4, 1, 1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, 3, 4, 4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, 3, 4, 4, 1, 1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, 3, 4, 4, 1, 1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, 3, 4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4, 3, 3, 4, 4, 1, 1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 Chlorophyll_WODflag =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 Chlorophyll_WODprofileflag = _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 Phaeophytin =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0.137, 0.129, 0.207, 0.236, 0.112, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _,
  0.137, 0.129, 0.207, 0.236, 0.112, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _,
  0.137, 0.129, 0.207, 0.236, 0.112, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _,
  0.137, 0.129, 0.207, 0.236, 0.112, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _,
  0.137, 0.129, 0.207, 0.236, 0.112, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _,
  0.137, 0.129, 0.207, 0.236, 0.112, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _,
  0.137, 0.129, 0.207, 0.236, 0.112, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _,
  0.137, 0.129, 0.207, 0.236, 0.112, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _,
  0.137, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  0.137, 0.129, 0.207, 0.236, 0.112, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _,
  0.137, 0.129, 0.207, 0.236, 0.112, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _,
  0.137, 0.129, 0.207, 0.236, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _,
  0.137, 0.129, 0.207, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _,
  0.137, 0.129, 0.207, 0.236, 0.112, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _,
  0.137, 0.129, 0.207, 0.236, 0.112, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _,
  0.271, 0.337, 0.5256667, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _,
  0.271, 0.337, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _,
  0.271, 0.337, 0.5256667, 0.236, 0.112, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _,
  0.271, 0.337, 0.5256667, 0.236, 0.112, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _,
  0.271, 0.337, 0.5256667, 0.236, 0.112, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _,
  0.271, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  0.271, 0.337, 0.5256667, 0.236, 0.112, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _,
  0.271, 0.337, 0.5256667, 0.236, 0.112, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _,
  0.271, 0.337, 0.5256667, 0.236, 0.112, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _,
  0.271, 0.337, 0.5256667, 0.236, 0.112, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _,
  0.271, 0.337, 0.5256667, 0.236, 0.112, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _,
  0.271, 0.337, 0.5256667, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _,
  0.271, 0.337, 0.5256667, 0.236, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _,
  0.271, 0.337, 0.5256667, 0.236, 0.112, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _,
  0.271, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  0.271, 0.337, 0.5256667, 0.236, 0.112, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _,
  0.271, 0.337, 0.5256667, 0.236, 0.112, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _,
  0.271, 0.337, 0.5256667, 0.236, 0.112, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _,
  0.271, 0.337, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _,
  0.271, 0.337, 0.5256667, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _,
  0.271, 0.337, 0.5256667, 0.236, 0.112, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _,
  0.271, 0.337, 0.5256667, 0.236, 0.112, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _,
  0.271, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  0.219, 0.137, 0.179, 0.216, 0.253, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _,
  0.219, 0.137, 0.179, 0.216, 0.253, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _,
  0.219, 0.137, 0.179, 0.216, 0.253, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _,
  0.219, 0.137, 0.179, 0.216, 0.253, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _,
  0.164, 0.082, 0.11, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _,
  0.164, 0.082, 0.11, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _,
  0.164, 0.082, 0.11, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _,
  0.164, 0.082, 0.11, 0.216, 0.253, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _,
  0.164, 0.082, 0.11, 0.216, 0.253, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _,
  0.164, 0.082, 0.11, 0.216, 0.253, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _,
  0.164, 0.082, 0.11, 0.216, 0.253, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _,
  0.164, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  0.164, 0.082, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _,
  0.164, 0.082, 0.11, 0.216, 0.253, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _,
  0.164, 0.082, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _,
  0.164, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  0.164, 0.082, 0.11, 0.216, 0.253, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _,
  0.164, 0.082, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _,
  0.164, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  0.164, 0.082, 0.11, 0.216, 0.253, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _,
  0.164, 0.082, 0.11, 0.216, 0.253, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _,
  0.164, 0.082, 0.11, 0.216, 0.253, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _,
  0.164, 0.082, 0.11, 0.216, 0.253, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _,
  0.164, 0.082, 0.11, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _,
  0.164, 0.082, 0.11, 0.216, 0.253, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _,
  0.344, 0.379, 0.3724074, 0.47, 0.898, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _,
  0.535, 0.31, 0.314, 0.191, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _,
  0.535, 0.31, 0.314, 0.191, 0.898, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _,
  0.535, 0.31, 0.314, 0.191, 0.898, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _,
  0.535, 0.31, 0.314, 0.191, 0.898, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _,
  0.535, 0.31, 0.314, 0.191, 0.898, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _,
  0.535, 0.31, 0.314, 0.191, 0.898, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _,
  0.535, 0.31, 0.314, 0.191, 0.898, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _,
  0.535, 0.31, 0.314, 0.191, 0.898, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _,
  0.535, 0.31, 0.314, 0.191, 0.898, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _,
  0.535, 0.31, 0.314, 0.191, 0.898, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _,
  0.535, 0.31, 0.314, 0.191, 0.898, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _,
  0.535, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  0.535, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  0.535, 0.31, 0.314, 0.191, 0.898, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _,
  0.535, 0.31, 0.314, 0.191, 0.898, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _,
  0.535, 0.31, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _,
  0.535, 0.31, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _,
  0.535, 0.31, 0.314, 0.191, 0.898, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _,
  0.535, 0.31, 0.314, 0.191, 0.898, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _,
  0.535, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  0.535, 0.31, 0.314, 0.191, 0.898, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _,
  0.535, 0.31, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _,
  0.535, 0.31, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _,
  0.535, 0.31, 0.314, 0.191, 0.898, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _,
  0.535, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  0.535, 0.31, 0.314, 0.191, 0.898, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _,
  0.535, 0.31, 0.314, 0.191, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _,
  0.535, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  0.392, 0.4, 0.361, 0.361, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _,
  0.392, 0.4, 0.361, 0.361, 0.898, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _,
  0.392, 0.4, 0.361, 0.361, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _,
  0.392, 0.4, 0.361, 0.361, 0.898, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _,
  0.392, 0.4, 0.361, 0.361, 0.898, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _,
  0.392, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  0.392, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  0.162, 0.113, 0.1665, 0.293, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _,
  0.162, 0.113, 0.1665, 0.293, 0.898, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _,
  0.162, 0.113, 0.1665, 0.293, 0.898, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _,
  0.162, 0.113, 0.1665, 0.293, 0.898, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _,
  0.162, 0.113, 0.1665, 0.293, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _,
  0.162, 0.113, 0.1665, 0.293, 0.898, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _,
  0.162, 0.113, 0.1665, 0.293, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _,
  0.162, 0.113, 0.1665, 0.293, 0.898, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _,
  0.162, 0.113, 0.1665, 0.293, 0.898, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _,
  0.162, 0.113, 0.1665, 0.293, 0.898, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _,
  0.162, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  0.253, 0.188, 0.18, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _,
  0.253, 0.188, 0.18, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _,
  0.253, 0.188, 0.18, 0.293, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _,
  0.253, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  0.253, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  0.253, 0.188, 0.18, 0.293, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _,
  0.253, 0.188, 0.18, 0.293, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _,
  0.253, 0.188, 0.18, 0.293, 0.898, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _,
  0.253, 0.188, 0.18, 0.293, 0.898, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _,
  0.253, 0.188, 0.18, 0.293, 0.898, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _,
  0.253, 0.188, 0.18, 0.293, 0.898, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _,
  0.253, 0.188, 0.18, 0.293, 0.898, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _,
  0.253, 0.188, 0.18, 0.293, 0.898, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _,
  0.253, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  0.253, 0.188, 0.18, 0.293, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _,
  0.253, 0.188, 0.18, 0.293, 0.898, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _,
  0.253, 0.188, 0.18, 0.293, 0.898, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _,
  0.253, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  0.094, 0.126, 0.141, 0.569, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _,
  0.094, 0.126, 0.141, 0.569, 0.898, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _,
  0.094, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  0.094, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  0.261, 0.327, 0.345, 0.354, 0.784, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _,
  0.261, 0.327, 0.345, 0.354, 0.784, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _,
  0.261, 0.327, 0.345, 0.354, 0.784, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _,
  0.261, 0.327, 0.345, 0.354, 0.784, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _,
  0.261, 0.327, 0.345, 0.354, 0.784, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _,
  0.261, 0.327, 0.345, 0.354, 0.784, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _,
  0.261, 0.327, 0.345, 0.354, 0.784, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _,
  0.261, 0.327, 0.345, 0.354, 0.784, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _,
  0.261, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  0.261, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  0.261, 0.327, 0.345, 0.354, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _,
  0.261, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  0.261, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  0.261, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  0.261, 0.327, 0.345, 0.354, 0.784, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _,
  0.261, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  0.261, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  0.261, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  0.261, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _ ;

 Phaeophytin_sigfigs =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, 3, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 Phaeophytin_WODflag =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 Alkalinity =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  2.238, 2.318, 2.337769, 2.340816, 2.349, 2.3515, 2.354, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _,
  2.238, 2.318, 2.337769, 2.340816, 2.349, 2.3515, 2.354, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _,
  2.238, 2.318, 2.337769, 2.340816, 2.349, 2.3515, 2.354, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _,
  2.238, 2.318, 2.337769, 2.340816, 2.349, 2.3515, 2.354, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _,
  2.238, 2.318, 2.337769, 2.340816, 2.349, 2.3515, 2.354, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _,
  2.238, 2.318, 2.337769, 2.340816, 2.349, 2.3515, 2.354, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _,
  2.238, 2.318, 2.337769, 2.340816, 2.349, 2.3515, 2.354, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _,
  2.238, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  2.238, 2.318, 2.337769, 2.340816, 2.349, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _,
  2.238, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  2.238, 2.318, 2.337769, 2.340816, 2.349, 2.3515, 2.354, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _,
  2.238, 2.318, 2.337769, 2.340816, 2.349, 2.3515, 2.354, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _,
  2.238, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  2.238, 2.318, 2.337769, 2.340816, 2.349, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _,
  2.238, 2.318, 2.337769, 2.340816, 2.349, 2.3515, 2.354, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _,
  2.238, 2.318, 2.337769, 2.340816, 2.349, 2.3515, 2.354, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _,
  2.238, 2.318, 2.337769, 2.340816, 2.349, 2.3515, 2.354, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _,
  2.238, 2.318, 2.337769, 2.340816, 2.349, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _,
  2.238, 2.318, 2.337769, 2.340816, 2.349, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _,
  2.238, 2.318, 2.337769, 2.340816, 2.349, 2.3515, 2.354, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _,
  2.238, 2.318, 2.337769, 2.340816, 2.349, 2.3515, 2.354, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _,
  2.238, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  2.238, 2.318, 2.337769, 2.340816, 2.349, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _,
  2.238, 2.318, 2.337769, 2.340816, 2.349, 2.3515, 2.354, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _,
  2.238, 2.318, 2.337769, 2.340816, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _,
  2.238, 2.318, 2.337769, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _,
  2.238, 2.318, 2.337769, 2.340816, 2.349, 2.3515, 2.354, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _,
  2.238, 2.318, 2.337769, 2.340816, 2.349, 2.3515, 2.354, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _,
  2.238, 2.318, 2.337769, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _,
  2.238, 2.318, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _,
  2.238, 2.318, 2.337769, 2.340816, 2.349, 2.3515, 2.354, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _,
  2.238, 2.318, 2.337769, 2.340816, 2.349, 2.3515, 2.354, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _,
  2.238, 2.318, 2.337769, 2.340816, 2.349, 2.3515, 2.354, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _,
  2.238, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  2.238, 2.318, 2.337769, 2.340816, 2.349, 2.3515, 2.354, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _,
  2.238, 2.318, 2.337769, 2.340816, 2.349, 2.3515, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _,
  2.238, 2.318, 2.337769, 2.340816, 2.349, 2.3515, 2.354, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _,
  2.238, 2.318, 2.337769, 2.340816, 2.349, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _,
  2.238, 2.318, 2.337769, 2.340816, 2.349, 2.3515, 2.354, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _,
  2.238, 2.318, 2.337769, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _,
  2.238, 2.318, 2.337769, 2.340816, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _,
  2.238, 2.318, 2.337769, 2.340816, 2.349, 2.3515, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _,
  2.238, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  2.238, 2.318, 2.337769, 2.340816, 2.349, 2.3515, 2.354, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _,
  2.238, 2.318, 2.337769, 2.340816, 2.349, 2.3515, 2.354, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _,
  2.238, 2.318, 2.337769, 2.340816, 2.349, 2.3515, 2.354, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _,
  2.238, 2.318, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _,
  2.238, 2.318, 2.337769, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _,
  2.238, 2.318, 2.337769, 2.340816, 2.349, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _,
  2.238, 2.318, 2.337769, 2.340816, 2.349, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _,
  2.238, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  2.238, 2.318, 2.337769, 2.340816, 2.349, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _,
  2.238, 2.318, 2.337769, 2.340816, 2.349, 2.3515, 2.354, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _,
  2.238, 2.318, 2.337769, 2.340816, 2.349, 2.3515, 2.354, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _,
  2.238, 2.318, 2.337769, 2.340816, 2.349, 2.3515, 2.354, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _,
  2.238, 2.318, 2.337769, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _,
  2.238, 2.318, 2.337769, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _,
  2.238, 2.318, 2.337769, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _,
  2.238, 2.318, 2.337769, 2.340816, 2.349, 2.3515, 2.354, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _,
  2.238, 2.318, 2.337769, 2.340816, 2.349, 2.3515, 2.354, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _,
  2.238, 2.318, 2.337769, 2.340816, 2.349, 2.3515, 2.354, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _,
  2.238, 2.318, 2.337769, 2.340816, 2.349, 2.3515, 2.354, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _,
  2.238, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  2.238, 2.318, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _,
  2.238, 2.318, 2.337769, 2.340816, 2.349, 2.3515, 2.354, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _,
  2.238, 2.318, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _,
  2.238, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  2.238, 2.318, 2.337769, 2.340816, 2.349, 2.3515, 2.354, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _,
  2.238, 2.318, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _,
  2.238, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  2.238, 2.318, 2.337769, 2.340816, 2.349, 2.3515, 2.354, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _,
  2.238, 2.318, 2.337769, 2.340816, 2.349, 2.3515, 2.354, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _,
  2.238, 2.318, 2.337769, 2.340816, 2.349, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _,
  2.238, 2.318, 2.337769, 2.340816, 2.349, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _,
  2.238, 2.318, 2.337769, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _,
  2.238, 2.318, 2.337769, 2.340816, 2.349, 2.3515, 2.354, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _,
  2.238, 2.318, 2.337769, 2.340816, 2.349, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _,
  2.238, 2.318, 2.337769, 2.340816, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _,
  2.238, 2.318, 2.337769, 2.340816, 2.349, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _,
  2.238, 2.318, 2.337769, 2.340816, 2.349, 2.3515, 2.354, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _,
  2.238, 2.318, 2.337769, 2.340816, 2.349, 2.3515, 2.354, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _,
  2.238, 2.318, 2.337769, 2.340816, 2.349, 2.3515, 2.354, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _,
  2.238, 2.318, 2.337769, 2.340816, 2.349, 2.3515, 2.354, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _,
  2.238, 2.318, 2.337769, 2.340816, 2.349, 2.3515, 2.354, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _,
  2.238, 2.318, 2.337769, 2.340816, 2.349, 2.3515, 2.354, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _,
  2.238, 2.318, 2.337769, 2.340816, 2.349, 2.3515, 2.354, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _,
  2.238, 2.318, 2.337769, 2.340816, 2.349, 2.3515, 2.354, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _,
  2.238, 2.318, 2.337769, 2.340816, 2.349, 2.3515, 2.354, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _,
  2.238, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  2.238, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  2.238, 2.318, 2.337769, 2.340816, 2.349, 2.3515, 2.354, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _,
  2.238, 2.318, 2.337769, 2.340816, 2.349, 2.3515, 2.354, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _,
  2.238, 2.318, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _,
  2.238, 2.318, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _,
  2.238, 2.318, 2.337769, 2.340816, 2.349, 2.3515, 2.354, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _,
  2.238, 2.318, 2.337769, 2.340816, 2.349, 2.3515, 2.354, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _,
  2.238, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  2.238, 2.318, 2.337769, 2.340816, 2.349, 2.3515, 2.354, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _,
  2.238, 2.318, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _,
  2.238, 2.318, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _,
  2.238, 2.318, 2.337769, 2.340816, 2.349, 2.3515, 2.354, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _,
  2.238, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  2.238, 2.318, 2.337769, 2.340816, 2.349, 2.3515, 2.354, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _,
  2.238, 2.318, 2.337769, 2.340816, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _,
  2.238, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  2.238, 2.318, 2.337769, 2.340816, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _,
  2.238, 2.318, 2.337769, 2.340816, 2.349, 2.3515, 2.354, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _,
  2.238, 2.318, 2.337769, 2.340816, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _,
  2.238, 2.318, 2.337769, 2.340816, 2.349, 2.3515, 2.354, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _,
  2.238, 2.318, 2.337769, 2.340816, 2.349, 2.3515, 2.354, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _,
  2.238, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  2.238, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  2.238, 2.318, 2.337769, 2.340816, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _,
  2.238, 2.318, 2.337769, 2.340816, 2.349, 2.3515, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _,
  2.238, 2.318, 2.337769, 2.340816, 2.349, 2.3515, 2.354, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _,
  2.238, 2.318, 2.337769, 2.340816, 2.349, 2.3515, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _,
  2.238, 2.318, 2.337769, 2.340816, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _,
  2.238, 2.318, 2.337769, 2.340816, 2.349, 2.3515, 2.354, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _,
  2.238, 2.318, 2.337769, 2.340816, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _,
  2.238, 2.318, 2.337769, 2.340816, 2.349, 2.3515, 2.354, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _,
  2.238, 2.318, 2.337769, 2.340816, 2.349, 2.3515, 2.354, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _,
  2.238, 2.318, 2.337769, 2.340816, 2.349, 2.3515, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _,
  2.238, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  2.238, 2.318, 2.337769, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _,
  2.238, 2.318, 2.337769, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _,
  2.238, 2.318, 2.337769, 2.340816, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _,
  2.238, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  2.238, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  2.238, 2.318, 2.337769, 2.340816, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _,
  2.238, 2.318, 2.337769, 2.340816, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _,
  2.238, 2.318, 2.337769, 2.340816, 2.349, 2.3515, 2.354, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _,
  2.238, 2.318, 2.337769, 2.340816, 2.349, 2.3515, 2.354, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _,
  2.238, 2.318, 2.337769, 2.340816, 2.349, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _,
  2.238, 2.318, 2.337769, 2.340816, 2.349, 2.3515, 2.354, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _,
  2.238, 2.318, 2.337769, 2.340816, 2.349, 2.3515, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _,
  2.238, 2.318, 2.337769, 2.340816, 2.349, 2.3515, 2.354, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _,
  2.238, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  2.238, 2.318, 2.337769, 2.340816, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _,
  2.238, 2.318, 2.337769, 2.340816, 2.349, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _,
  2.238, 2.318, 2.337769, 2.340816, 2.349, 2.3515, 2.354, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _,
  2.238, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  2.238, 2.318, 2.337769, 2.340816, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _,
  2.238, 2.318, 2.337769, 2.340816, 2.349, 2.3515, 2.354, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _,
  2.238, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  2.238, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  2.238, 2.318, 2.337769, 2.340816, 2.349, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _,
  2.238, 2.318, 2.337769, 2.340816, 2.349, 2.3515, 2.354, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _,
  2.238, 2.318, 2.337769, 2.340816, 2.349, 2.3515, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _,
  2.238, 2.318, 2.337769, 2.340816, 2.349, 2.3515, 2.354, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _,
  2.238, 2.318, 2.337769, 2.340816, 2.349, 2.3515, 2.354, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _,
  2.238, 2.318, 2.337769, 2.340816, 2.349, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _,
  2.238, 2.318, 2.337769, 2.340816, 2.349, 2.3515, 2.354, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _,
  2.238, 2.318, 2.337769, 2.340816, 2.349, 2.3515, 2.354, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _,
  2.238, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  2.238, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  2.238, 2.318, 2.337769, 2.340816, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _,
  2.238, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  2.238, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  2.238, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  2.238, 2.318, 2.337769, 2.340816, 2.349, 2.3515, 2.354, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _,
  2.238, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  2.238, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  2.238, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  2.238, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _ ;

 Alkalinity_sigfigs =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4, 4, 4, 4, 4, 4, 4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4, 4, 4, 4, 4, 4, 4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4, 4, 4, 4, 4, 4, 4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4, 4, 4, 4, 4, 4, 4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4, 4, 4, 4, 4, 4, 4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4, 4, 4, 4, 4, 4, 4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4, 4, 4, 4, 4, 4, 4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4, 4, 4, 4, 4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4, 4, 4, 4, 4, 4, 4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4, 4, 4, 4, 4, 4, 4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4, 4, 4, 4, 4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4, 4, 4, 4, 4, 4, 4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4, 4, 4, 4, 4, 4, 4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4, 4, 4, 4, 4, 4, 4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4, 4, 4, 4, 4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4, 4, 4, 4, 4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4, 4, 4, 4, 4, 4, 4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4, 4, 4, 4, 4, 4, 4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4, 4, 4, 4, 4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4, 4, 4, 4, 4, 4, 4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4, 4, 4, 4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4, 4, 4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4, 4, 4, 4, 4, 4, 4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4, 4, 4, 4, 4, 4, 4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4, 4, 4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4, 4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4, 4, 4, 4, 4, 4, 4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4, 4, 4, 4, 4, 4, 4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4, 4, 4, 4, 4, 4, 4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4, 4, 4, 4, 4, 4, 4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4, 4, 4, 4, 4, 4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4, 4, 4, 4, 4, 4, 4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4, 4, 4, 4, 4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4, 4, 4, 4, 4, 4, 4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4, 4, 4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4, 4, 4, 4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4, 4, 4, 4, 4, 4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4, 4, 4, 4, 4, 4, 4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4, 4, 4, 4, 4, 4, 4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4, 4, 4, 4, 4, 4, 4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4, 4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4, 4, 4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4, 4, 4, 4, 4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4, 4, 4, 4, 4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4, 4, 4, 4, 4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4, 4, 4, 4, 4, 4, 4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4, 4, 4, 4, 4, 4, 4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4, 4, 4, 4, 4, 4, 4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4, 4, 4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4, 4, 4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4, 4, 4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4, 4, 4, 4, 4, 4, 4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4, 4, 4, 4, 4, 4, 4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4, 4, 4, 4, 4, 4, 4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4, 4, 4, 4, 4, 4, 4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4, 4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4, 4, 4, 4, 4, 4, 4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4, 4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4, 4, 4, 4, 4, 4, 4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4, 4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4, 4, 4, 4, 4, 4, 4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4, 4, 4, 4, 4, 4, 4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4, 4, 4, 4, 4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4, 4, 4, 4, 4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4, 4, 4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4, 4, 4, 4, 4, 4, 4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4, 4, 4, 4, 4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4, 4, 4, 4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4, 4, 4, 4, 4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4, 4, 4, 4, 4, 4, 4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4, 4, 4, 4, 4, 4, 4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4, 4, 4, 4, 4, 4, 4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4, 4, 4, 4, 4, 4, 4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4, 4, 4, 4, 4, 4, 4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4, 4, 4, 4, 4, 4, 4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4, 4, 4, 4, 4, 4, 4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4, 4, 4, 4, 4, 4, 4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4, 4, 4, 4, 4, 4, 4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4, 4, 4, 4, 4, 4, 4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4, 4, 4, 4, 4, 4, 4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4, 4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4, 4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4, 4, 4, 4, 4, 4, 4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4, 4, 4, 4, 4, 4, 4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4, 4, 4, 4, 4, 4, 4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4, 4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4, 4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4, 4, 4, 4, 4, 4, 4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4, 4, 4, 4, 4, 4, 4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4, 4, 4, 4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4, 4, 4, 4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4, 4, 4, 4, 4, 4, 4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4, 4, 4, 4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4, 4, 4, 4, 4, 4, 4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4, 4, 4, 4, 4, 4, 4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4, 4, 4, 4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4, 4, 4, 4, 4, 4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4, 4, 4, 4, 4, 4, 4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4, 4, 4, 4, 4, 4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4, 4, 4, 4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4, 4, 4, 4, 4, 4, 4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4, 4, 4, 4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4, 4, 4, 4, 4, 4, 4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4, 4, 4, 4, 4, 4, 4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4, 4, 4, 4, 4, 4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4, 4, 4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4, 4, 4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4, 4, 4, 4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4, 4, 4, 4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4, 4, 4, 4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4, 4, 4, 4, 4, 4, 4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4, 4, 4, 4, 4, 4, 4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4, 4, 4, 4, 4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4, 4, 4, 4, 4, 4, 4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4, 4, 4, 4, 4, 4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4, 4, 4, 4, 4, 4, 4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4, 4, 4, 4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4, 4, 4, 4, 4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4, 4, 4, 4, 4, 4, 4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4, 4, 4, 4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4, 4, 4, 4, 4, 4, 4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4, 4, 4, 4, 4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4, 4, 4, 4, 4, 4, 4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4, 4, 4, 4, 4, 4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4, 4, 4, 4, 4, 4, 4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4, 4, 4, 4, 4, 4, 4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4, 4, 4, 4, 4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4, 4, 4, 4, 4, 4, 4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4, 4, 4, 4, 4, 4, 4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4, 4, 4, 4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4, 4, 4, 4, 4, 4, 4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 Alkalinity_WODflag =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 Alkalinity_WODprofileflag = _, _, _, _, _, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 NO2NO3 =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 0.18, 0.15, 0.86, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _,
  _, 0.18, 0.15, 0.86, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _,
  _, 0.18, 0.15, 0.86, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _,
  _, 0.18, 0.15, 0.86, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _,
  _, 0.18, 0.15, 0.86, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _,
  _, 0.18, 0.15, 0.86, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _,
  _, 0.18, 0.15, 0.86, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _,
  _, 0.18, 0.15, 0.86, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 0.18, 0.15, 0.86, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 0.18, 0.15, 0.86, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _,
  _, 0.18, 0.15, 0.86, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 0.18, 0.15, 0.86, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _,
  _, 0.18, 0.15, 0.86, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _,
  _, 0.18, 0.15, 0.86, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _,
  _, 0.18, 0.15, 0.86, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _,
  _, 0.18, 0.15, 0.86, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _,
  _, 0.18, 0.15, 0.86, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _,
  _, 0.18, 0.15, 0.86, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _,
  _, 0.18, 0.15, 0.86, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 0.18, 0.15, 0.86, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _,
  _, 0.18, 0.15, 0.86, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _,
  _, 0.18, 0.15, 0.86, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _,
  _, 0.18, 0.15, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _,
  _, 0.18, 0.15, 0.86, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _,
  _, 0.18, 0.15, 0.86, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _,
  _, 0.18, 0.15, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _,
  _, 0.18, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  _, 0.18, 0.15, 0.86, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _,
  _, 0.18, 0.15, 0.86, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _,
  _, 0.18, 0.15, 0.86, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 0.18, 0.15, 0.86, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _,
  _, 0.18, 0.15, 0.86, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _,
  _, 0.18, 0.15, 0.86, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _,
  _, 0.18, 0.15, 0.86, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _,
  _, 0.18, 0.15, 0.86, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _,
  _, 0.18, 0.15, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _,
  _, 0.18, 0.15, 0.86, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _,
  _, 0.18, 0.15, 0.86, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 0.18, 0.15, 0.86, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _,
  _, 0.18, 0.15, 0.86, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _,
  _, 0.18, 0.15, 0.86, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _,
  _, 0.18, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  _, 0.18, 0.15, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _,
  _, 0.18, 0.15, 0.86, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _,
  _, 0.18, 0.15, 0.86, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 0.18, 0.15, 0.86, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _,
  _, 0.18, 0.15, 0.86, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _,
  _, 0.18, 0.15, 0.86, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _,
  _, 0.18, 0.15, 0.86, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _,
  _, 0.18, 0.15, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _,
  _, 0.18, 0.15, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _,
  _, 0.18, 0.15, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _,
  _, 0.18, 0.15, 0.86, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _,
  _, 0.18, 0.15, 0.86, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _,
  _, 0.18, 0.15, 0.86, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _,
  _, 0.18, 0.15, 0.86, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 0.18, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  _, 0.18, 0.15, 0.86, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _,
  _, 0.18, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 0.18, 0.15, 0.86, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _,
  _, 0.18, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 0.18, 0.15, 0.86, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _,
  _, 0.18, 0.15, 0.86, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _,
  _, 0.18, 0.15, 0.86, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _,
  _, 0.18, 0.15, 0.86, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _,
  _, 0.18, 0.15, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _,
  _, 0.18, 0.15, 0.86, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _,
  _, 0.18, 0.15, 0.86, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _,
  _, 0.18, 0.15, 0.86, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _,
  _, 0.18, 0.15, 0.86, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _,
  _, 0.18, 0.15, 0.86, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _,
  _, 0.18, 0.15, 0.86, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _,
  _, 0.18, 0.15, 0.86, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _,
  _, 0.18, 0.15, 0.86, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _,
  _, 0.18, 0.15, 0.86, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _,
  _, 0.18, 0.15, 0.86, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _,
  _, 0.18, 0.15, 0.86, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _,
  _, 0.18, 0.15, 0.86, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _,
  _, 0.18, 0.15, 0.86, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 0.18, 0.15, 0.86, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _,
  _, 0.18, 0.15, 0.86, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _,
  _, 0.18, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  _, 0.18, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  _, 0.18, 0.15, 0.86, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _,
  _, 0.18, 0.15, 0.86, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 0.18, 0.15, 0.86, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _,
  _, 0.18, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  _, 0.18, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  _, 0.18, 0.15, 0.86, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 0.18, 0.15, 0.86, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _,
  _, 0.18, 0.15, 0.86, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 0.18, 0.15, 0.86, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _,
  _, 0.18, 0.15, 0.86, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _,
  _, 0.18, 0.15, 0.86, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _,
  _, 0.18, 0.15, 0.86, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _,
  _, 0.18, 0.15, 0.86, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 0.18, 0.15, 0.86, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _,
  _, 0.18, 0.15, 0.86, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _,
  _, 0.18, 0.15, 0.86, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _,
  _, 0.18, 0.15, 0.86, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _,
  _, 0.18, 0.15, 0.86, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _,
  _, 0.18, 0.15, 0.86, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _,
  _, 0.18, 0.15, 0.86, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _,
  _, 0.18, 0.15, 0.86, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _,
  _, 0.18, 0.15, 0.86, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _,
  _, 0.18, 0.15, 0.86, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 0.18, 0.15, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _,
  _, 0.18, 0.15, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _,
  _, 0.18, 0.15, 0.86, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 0.18, 0.15, 0.86, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _,
  _, 0.18, 0.15, 0.86, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _,
  _, 0.18, 0.15, 0.86, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _,
  _, 0.18, 0.15, 0.86, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _,
  _, 0.18, 0.15, 0.86, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _,
  _, 0.18, 0.15, 0.86, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _,
  _, 0.18, 0.15, 0.86, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _,
  _, 0.18, 0.15, 0.86, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 0.18, 0.15, 0.86, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _,
  _, 0.18, 0.15, 0.86, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _,
  _, 0.18, 0.15, 0.86, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 0.18, 0.15, 0.86, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _,
  _, 0.18, 0.15, 0.86, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 0.18, 0.15, 0.86, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _,
  _, 0.18, 0.15, 0.86, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _,
  _, 0.18, 0.15, 0.86, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _,
  _, 0.18, 0.15, 0.86, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _,
  _, 0.18, 0.15, 0.86, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _,
  _, 0.18, 0.15, 0.86, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _,
  _, 0.18, 0.15, 0.86, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _,
  _, 0.18, 0.15, 0.86, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 0.18, 0.15, 0.86, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 0.18, 0.15, 0.86, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 NO2NO3_sigfigs =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 3, 3, 3, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 NO2NO3_WODflag =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 crs = _ ;

 WODf = _ ;

 WODfp = _ ;

 WODfd = _ ;
}

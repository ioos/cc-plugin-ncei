netcdf Kachemak_Bay { 
dimensions:
   Sample_Site = 34 ;
   NST_Site_code_string_length = 8 ;
   Site_name_string_length = 30 ;
variables:
   double Ampelisca_Survival___mean(Sample_Site) ;
      Ampelisca_Survival___mean:long_name = "Ampelisca Survival - mean" ;
      Ampelisca_Survival___mean:coordinates = "latitude longitude time z" ;
      Ampelisca_Survival___mean:matix = "SED" ;
      Ampelisca_Survival___mean:units = "percent" ;
      Ampelisca_Survival___mean:_FillValue = -1. ;
      Ampelisca_Survival___mean:valid_min = 0. ;
      Ampelisca_Survival___mean:valid_max = 100. ;
      Ampelisca_Survival___mean:instrument = "AMP_AA" ;
      Ampelisca_Survival___mean:grid_mapping = "crs" ;
      Ampelisca_Survival___mean:reference = "0074376/data/0-data/Bioeffects_Assessments/Kachemak_Bay/Data_Files/KB1_ASSAY.txt" ;
   double Ampelisca_Survival___standard_deviation(Sample_Site) ;
      Ampelisca_Survival___standard_deviation:long_name = "Ampelisca Survival - standard deviation" ;
      Ampelisca_Survival___standard_deviation:coordinates = "latitude longitude time z" ;
      Ampelisca_Survival___standard_deviation:matix = "SED" ;
      Ampelisca_Survival___standard_deviation:units = "count/count" ;
      Ampelisca_Survival___standard_deviation:_FillValue = -1. ;
      Ampelisca_Survival___standard_deviation:valid_min = 0. ;
      Ampelisca_Survival___standard_deviation:valid_max = 1.79769313486232e+308 ;
      Ampelisca_Survival___standard_deviation:instrument = "AMP_AA" ;
      Ampelisca_Survival___standard_deviation:grid_mapping = "crs" ;
      Ampelisca_Survival___standard_deviation:reference = "0074376/data/0-data/Bioeffects_Assessments/Kachemak_Bay/Data_Files/KB1_ASSAY.txt" ;
   double Ampelisca_Survival_as___of_Control___mean(Sample_Site) ;
      Ampelisca_Survival_as___of_Control___mean:long_name = "Ampelisca Survival as % of Control - mean" ;
      Ampelisca_Survival_as___of_Control___mean:coordinates = "latitude longitude time z" ;
      Ampelisca_Survival_as___of_Control___mean:matix = "SED" ;
      Ampelisca_Survival_as___of_Control___mean:units = "percent" ;
      Ampelisca_Survival_as___of_Control___mean:_FillValue = -1. ;
      Ampelisca_Survival_as___of_Control___mean:valid_min = 0. ;
      Ampelisca_Survival_as___of_Control___mean:valid_max = 100. ;
      Ampelisca_Survival_as___of_Control___mean:instrument = "AMP_AA" ;
      Ampelisca_Survival_as___of_Control___mean:grid_mapping = "crs" ;
      Ampelisca_Survival_as___of_Control___mean:reference = "0074376/data/0-data/Bioeffects_Assessments/Kachemak_Bay/Data_Files/KB1_ASSAY.txt" ;
   double Eohaustorius_Survival___standard_deviation(Sample_Site) ;
      Eohaustorius_Survival___standard_deviation:long_name = "Eohaustorius Survival - standard deviation" ;
      Eohaustorius_Survival___standard_deviation:coordinates = "latitude longitude time z" ;
      Eohaustorius_Survival___standard_deviation:matix = "SED" ;
      Eohaustorius_Survival___standard_deviation:units = "count/count" ;
      Eohaustorius_Survival___standard_deviation:_FillValue = -1. ;
      Eohaustorius_Survival___standard_deviation:valid_min = 0. ;
      Eohaustorius_Survival___standard_deviation:valid_max = 1.79769313486232e+308 ;
      Eohaustorius_Survival___standard_deviation:instrument = "AMP_EE" ;
      Eohaustorius_Survival___standard_deviation:grid_mapping = "crs" ;
      Eohaustorius_Survival___standard_deviation:reference = "0074376/data/0-data/Bioeffects_Assessments/Kachemak_Bay/Data_Files/KB1_ASSAY.txt" ;
   double Eohaustorius_mean_survival(Sample_Site) ;
      Eohaustorius_mean_survival:long_name = "Eohaustorius mean survival" ;
      Eohaustorius_mean_survival:coordinates = "latitude longitude time z" ;
      Eohaustorius_mean_survival:matix = "SED" ;
      Eohaustorius_mean_survival:units = "percent" ;
      Eohaustorius_mean_survival:_FillValue = -1. ;
      Eohaustorius_mean_survival:valid_min = 0. ;
      Eohaustorius_mean_survival:valid_max = 100. ;
      Eohaustorius_mean_survival:instrument = "AMP_EE" ;
      Eohaustorius_mean_survival:grid_mapping = "crs" ;
      Eohaustorius_mean_survival:reference = "0074376/data/0-data/Bioeffects_Assessments/Kachemak_Bay/Data_Files/KB1_ASSAY.txt" ;
   double Eohaustorius_survival_count(Sample_Site) ;
      Eohaustorius_survival_count:long_name = "Eohaustorius survival count" ;
      Eohaustorius_survival_count:coordinates = "latitude longitude time z" ;
      Eohaustorius_survival_count:matix = "SED" ;
      Eohaustorius_survival_count:units = "count" ;
      Eohaustorius_survival_count:_FillValue = -1. ;
      Eohaustorius_survival_count:valid_min = 0. ;
      Eohaustorius_survival_count:valid_max = 1.79769313486232e+308 ;
      Eohaustorius_survival_count:instrument = "AMP_EE" ;
      Eohaustorius_survival_count:grid_mapping = "crs" ;
      Eohaustorius_survival_count:reference = "0074376/data/0-data/Bioeffects_Assessments/Kachemak_Bay/Data_Files/KB1_ASSAY.txt" ;
   double Density___mean(Sample_Site) ;
      Density___mean:long_name = "Density - mean" ;
      Density___mean:coordinates = "latitude longitude time z" ;
      Density___mean:matix = "SED" ;
      Density___mean:units = "count" ;
      Density___mean:_FillValue = -1. ;
      Density___mean:valid_min = 0. ;
      Density___mean:valid_max = 1.79769313486232e+308 ;
      Density___mean:instrument = "" ;
      Density___mean:grid_mapping = "crs" ;
      Density___mean:reference = "0074376/data/0-data/Bioeffects_Assessments/Kachemak_Bay/Data_Files/KB1_BENTHIC.txt" ;
   double Diversity(Sample_Site) ;
      Diversity:long_name = "Diversity" ;
      Diversity:coordinates = "latitude longitude time z" ;
      Diversity:matix = "SED" ;
      Diversity:units = "count" ;
      Diversity:_FillValue = -1. ;
      Diversity:valid_min = 0. ;
      Diversity:valid_max = 1.79769313486232e+308 ;
      Diversity:instrument = "" ;
      Diversity:grid_mapping = "crs" ;
      Diversity:reference = "0074376/data/0-data/Bioeffects_Assessments/Kachemak_Bay/Data_Files/KB1_BENTHIC.txt" ;
   double Evenness(Sample_Site) ;
      Evenness:long_name = "Evenness" ;
      Evenness:coordinates = "latitude longitude time z" ;
      Evenness:matix = "SED" ;
      Evenness:units = "count" ;
      Evenness:_FillValue = -1. ;
      Evenness:valid_min = 0. ;
      Evenness:valid_max = 1.79769313486232e+308 ;
      Evenness:instrument = "" ;
      Evenness:grid_mapping = "crs" ;
      Evenness:reference = "0074376/data/0-data/Bioeffects_Assessments/Kachemak_Bay/Data_Files/KB1_BENTHIC.txt" ;
   double Individuals___total(Sample_Site) ;
      Individuals___total:long_name = "Individuals - total" ;
      Individuals___total:coordinates = "latitude longitude time z" ;
      Individuals___total:matix = "SED" ;
      Individuals___total:units = "count" ;
      Individuals___total:_FillValue = -1. ;
      Individuals___total:valid_min = 0. ;
      Individuals___total:valid_max = 1.79769313486232e+308 ;
      Individuals___total:instrument = "" ;
      Individuals___total:grid_mapping = "crs" ;
      Individuals___total:reference = "0074376/data/0-data/Bioeffects_Assessments/Kachemak_Bay/Data_Files/KB1_BENTHIC.txt" ;
   double Taxa___Total(Sample_Site) ;
      Taxa___Total:long_name = "Taxa - Total" ;
      Taxa___Total:coordinates = "latitude longitude time z" ;
      Taxa___Total:matix = "SED" ;
      Taxa___Total:units = "count" ;
      Taxa___Total:_FillValue = -1. ;
      Taxa___Total:valid_min = 0. ;
      Taxa___Total:valid_max = 1.79769313486232e+308 ;
      Taxa___Total:instrument = "" ;
      Taxa___Total:grid_mapping = "crs" ;
      Taxa___Total:reference = "0074376/data/0-data/Bioeffects_Assessments/Kachemak_Bay/Data_Files/KB1_BENTHIC.txt" ;
   double Clostridium_perfringens___dry(Sample_Site) ;
      Clostridium_perfringens___dry:long_name = "Clostridium perfringens - dry" ;
      Clostridium_perfringens___dry:coordinates = "latitude longitude time z" ;
      Clostridium_perfringens___dry:matix = "SED" ;
      Clostridium_perfringens___dry:units = "count/gram" ;
      Clostridium_perfringens___dry:_FillValue = -1. ;
      Clostridium_perfringens___dry:valid_min = 0. ;
      Clostridium_perfringens___dry:valid_max = 1.79769313486232e+308 ;
      Clostridium_perfringens___dry:instrument = "" ;
      Clostridium_perfringens___dry:grid_mapping = "crs" ;
      Clostridium_perfringens___dry:reference = "0074376/data/0-data/Bioeffects_Assessments/Kachemak_Bay/Data_Files/KB1_C_PERF.txt" ;
   double Clostridium_perfringens___wet(Sample_Site) ;
      Clostridium_perfringens___wet:long_name = "Clostridium perfringens - wet" ;
      Clostridium_perfringens___wet:coordinates = "latitude longitude time z" ;
      Clostridium_perfringens___wet:matix = "SED" ;
      Clostridium_perfringens___wet:units = "count/gram" ;
      Clostridium_perfringens___wet:_FillValue = -1. ;
      Clostridium_perfringens___wet:valid_min = 0. ;
      Clostridium_perfringens___wet:valid_max = 1.79769313486232e+308 ;
      Clostridium_perfringens___wet:instrument = "" ;
      Clostridium_perfringens___wet:grid_mapping = "crs" ;
      Clostridium_perfringens___wet:reference = "0074376/data/0-data/Bioeffects_Assessments/Kachemak_Bay/Data_Files/KB1_C_PERF.txt" ;
   double Clostridium_perfrirgens___Count_1(Sample_Site) ;
      Clostridium_perfrirgens___Count_1:long_name = "Clostridium perfrirgens - Count 1" ;
      Clostridium_perfrirgens___Count_1:coordinates = "latitude longitude time z" ;
      Clostridium_perfrirgens___Count_1:matix = "SED" ;
      Clostridium_perfrirgens___Count_1:units = "count" ;
      Clostridium_perfrirgens___Count_1:_FillValue = -1. ;
      Clostridium_perfrirgens___Count_1:valid_min = 0. ;
      Clostridium_perfrirgens___Count_1:valid_max = 1.79769313486232e+308 ;
      Clostridium_perfrirgens___Count_1:instrument = "" ;
      Clostridium_perfrirgens___Count_1:grid_mapping = "crs" ;
      Clostridium_perfrirgens___Count_1:reference = "0074376/data/0-data/Bioeffects_Assessments/Kachemak_Bay/Data_Files/KB1_C_PERF.txt" ;
   double Clostridium_perfrirgens___Count_2(Sample_Site) ;
      Clostridium_perfrirgens___Count_2:long_name = "Clostridium perfrirgens - Count 2" ;
      Clostridium_perfrirgens___Count_2:coordinates = "latitude longitude time z" ;
      Clostridium_perfrirgens___Count_2:matix = "SED" ;
      Clostridium_perfrirgens___Count_2:units = "count" ;
      Clostridium_perfrirgens___Count_2:_FillValue = -1. ;
      Clostridium_perfrirgens___Count_2:valid_min = 0. ;
      Clostridium_perfrirgens___Count_2:valid_max = 1.79769313486232e+308 ;
      Clostridium_perfrirgens___Count_2:instrument = "" ;
      Clostridium_perfrirgens___Count_2:grid_mapping = "crs" ;
      Clostridium_perfrirgens___Count_2:reference = "0074376/data/0-data/Bioeffects_Assessments/Kachemak_Bay/Data_Files/KB1_C_PERF.txt" ;
   double Clostridium_perfrirgens___Mean(Sample_Site) ;
      Clostridium_perfrirgens___Mean:long_name = "Clostridium perfrirgens - Mean" ;
      Clostridium_perfrirgens___Mean:coordinates = "latitude longitude time z" ;
      Clostridium_perfrirgens___Mean:matix = "SED" ;
      Clostridium_perfrirgens___Mean:units = "count" ;
      Clostridium_perfrirgens___Mean:_FillValue = -1. ;
      Clostridium_perfrirgens___Mean:valid_min = 0. ;
      Clostridium_perfrirgens___Mean:valid_max = 1.79769313486232e+308 ;
      Clostridium_perfrirgens___Mean:instrument = "" ;
      Clostridium_perfrirgens___Mean:grid_mapping = "crs" ;
      Clostridium_perfrirgens___Mean:reference = "0074376/data/0-data/Bioeffects_Assessments/Kachemak_Bay/Data_Files/KB1_C_PERF.txt" ;
   double Clostridium_perfrirgens___Moisture(Sample_Site) ;
      Clostridium_perfrirgens___Moisture:long_name = "Clostridium perfrirgens - Moisture" ;
      Clostridium_perfrirgens___Moisture:coordinates = "latitude longitude time z" ;
      Clostridium_perfrirgens___Moisture:matix = "SED" ;
      Clostridium_perfrirgens___Moisture:units = "percent" ;
      Clostridium_perfrirgens___Moisture:_FillValue = -1. ;
      Clostridium_perfrirgens___Moisture:valid_min = 0. ;
      Clostridium_perfrirgens___Moisture:valid_max = 100. ;
      Clostridium_perfrirgens___Moisture:instrument = "" ;
      Clostridium_perfrirgens___Moisture:grid_mapping = "crs" ;
      Clostridium_perfrirgens___Moisture:reference = "0074376/data/0-data/Bioeffects_Assessments/Kachemak_Bay/Data_Files/KB1_C_PERF.txt" ;
   double Chemical_1_2_3_4_Tetrachlorobenzene(Sample_Site) ;
      Chemical_1_2_3_4_Tetrachlorobenzene:long_name = "1,2,3,4-Tetrachlorobenzene" ;
      Chemical_1_2_3_4_Tetrachlorobenzene:coordinates = "latitude longitude time z" ;
      Chemical_1_2_3_4_Tetrachlorobenzene:matix = "SED" ;
      Chemical_1_2_3_4_Tetrachlorobenzene:units = "nanograms/gram" ;
      Chemical_1_2_3_4_Tetrachlorobenzene:_FillValue = -1. ;
      Chemical_1_2_3_4_Tetrachlorobenzene:valid_min = 0. ;
      Chemical_1_2_3_4_Tetrachlorobenzene:valid_max = 1.79769313486232e+308 ;
      Chemical_1_2_3_4_Tetrachlorobenzene:instrument = "ECDDUAL_M_Sample_dry_weight" ;
      Chemical_1_2_3_4_Tetrachlorobenzene:grid_mapping = "crs" ;
      Chemical_1_2_3_4_Tetrachlorobenzene:reference = "0074376/data/0-data/Bioeffects_Assessments/Kachemak_Bay/Data_Files/KB1_ORG.txt" ;
   double Chemical_1_2_4_5_Tetrachlorobenzene(Sample_Site) ;
      Chemical_1_2_4_5_Tetrachlorobenzene:long_name = "1,2,4,5-Tetrachlorobenzene" ;
      Chemical_1_2_4_5_Tetrachlorobenzene:coordinates = "latitude longitude time z" ;
      Chemical_1_2_4_5_Tetrachlorobenzene:matix = "SED" ;
      Chemical_1_2_4_5_Tetrachlorobenzene:units = "nanograms/gram" ;
      Chemical_1_2_4_5_Tetrachlorobenzene:_FillValue = -1. ;
      Chemical_1_2_4_5_Tetrachlorobenzene:valid_min = 0. ;
      Chemical_1_2_4_5_Tetrachlorobenzene:valid_max = 1.79769313486232e+308 ;
      Chemical_1_2_4_5_Tetrachlorobenzene:instrument = "ECDDUAL_M_Sample_dry_weight" ;
      Chemical_1_2_4_5_Tetrachlorobenzene:grid_mapping = "crs" ;
      Chemical_1_2_4_5_Tetrachlorobenzene:reference = "0074376/data/0-data/Bioeffects_Assessments/Kachemak_Bay/Data_Files/KB1_ORG.txt" ;
   double Chemical_2_4__DDD(Sample_Site) ;
      Chemical_2_4__DDD:long_name = "2,4\'-DDD" ;
      Chemical_2_4__DDD:coordinates = "latitude longitude time z" ;
      Chemical_2_4__DDD:matix = "SED" ;
      Chemical_2_4__DDD:units = "nanograms/gram" ;
      Chemical_2_4__DDD:_FillValue = -1. ;
      Chemical_2_4__DDD:valid_min = 0. ;
      Chemical_2_4__DDD:valid_max = 1.79769313486232e+308 ;
      Chemical_2_4__DDD:instrument = "ECDDUAL_M_Sample_dry_weight" ;
      Chemical_2_4__DDD:grid_mapping = "crs" ;
      Chemical_2_4__DDD:reference = "0074376/data/0-data/Bioeffects_Assessments/Kachemak_Bay/Data_Files/KB1_ORG.txt" ;
   double Chemical_2_4__DDE(Sample_Site) ;
      Chemical_2_4__DDE:long_name = "2,4\'-DDE" ;
      Chemical_2_4__DDE:coordinates = "latitude longitude time z" ;
      Chemical_2_4__DDE:matix = "SED" ;
      Chemical_2_4__DDE:units = "nanograms/gram" ;
      Chemical_2_4__DDE:_FillValue = -1. ;
      Chemical_2_4__DDE:valid_min = 0. ;
      Chemical_2_4__DDE:valid_max = 1.79769313486232e+308 ;
      Chemical_2_4__DDE:instrument = "ECDDUAL_M_Sample_dry_weight" ;
      Chemical_2_4__DDE:grid_mapping = "crs" ;
      Chemical_2_4__DDE:reference = "0074376/data/0-data/Bioeffects_Assessments/Kachemak_Bay/Data_Files/KB1_ORG.txt" ;
   double Chemical_2_4__DDT(Sample_Site) ;
      Chemical_2_4__DDT:long_name = "2,4\'-DDT" ;
      Chemical_2_4__DDT:coordinates = "latitude longitude time z" ;
      Chemical_2_4__DDT:matix = "SED" ;
      Chemical_2_4__DDT:units = "nanograms/gram" ;
      Chemical_2_4__DDT:_FillValue = -1. ;
      Chemical_2_4__DDT:valid_min = 0. ;
      Chemical_2_4__DDT:valid_max = 1.79769313486232e+308 ;
      Chemical_2_4__DDT:instrument = "ECDDUAL_M_Sample_dry_weight" ;
      Chemical_2_4__DDT:grid_mapping = "crs" ;
      Chemical_2_4__DDT:reference = "0074376/data/0-data/Bioeffects_Assessments/Kachemak_Bay/Data_Files/KB1_ORG.txt" ;
   double Chemical_4_4__DDD(Sample_Site) ;
      Chemical_4_4__DDD:long_name = "4,4\'-DDD" ;
      Chemical_4_4__DDD:coordinates = "latitude longitude time z" ;
      Chemical_4_4__DDD:matix = "SED" ;
      Chemical_4_4__DDD:units = "nanograms/gram" ;
      Chemical_4_4__DDD:_FillValue = -1. ;
      Chemical_4_4__DDD:valid_min = 0. ;
      Chemical_4_4__DDD:valid_max = 1.79769313486232e+308 ;
      Chemical_4_4__DDD:instrument = "ECDDUAL_M_Sample_dry_weight" ;
      Chemical_4_4__DDD:grid_mapping = "crs" ;
      Chemical_4_4__DDD:reference = "0074376/data/0-data/Bioeffects_Assessments/Kachemak_Bay/Data_Files/KB1_ORG.txt" ;
   double Chemical_4_4__DDE(Sample_Site) ;
      Chemical_4_4__DDE:long_name = "4,4\'-DDE" ;
      Chemical_4_4__DDE:coordinates = "latitude longitude time z" ;
      Chemical_4_4__DDE:matix = "SED" ;
      Chemical_4_4__DDE:units = "nanograms/gram" ;
      Chemical_4_4__DDE:_FillValue = -1. ;
      Chemical_4_4__DDE:valid_min = 0. ;
      Chemical_4_4__DDE:valid_max = 1.79769313486232e+308 ;
      Chemical_4_4__DDE:instrument = "ECDDUAL_M_Sample_dry_weight" ;
      Chemical_4_4__DDE:grid_mapping = "crs" ;
      Chemical_4_4__DDE:reference = "0074376/data/0-data/Bioeffects_Assessments/Kachemak_Bay/Data_Files/KB1_ORG.txt" ;
   double Chemical_4_4__DDT(Sample_Site) ;
      Chemical_4_4__DDT:long_name = "4,4\'-DDT" ;
      Chemical_4_4__DDT:coordinates = "latitude longitude time z" ;
      Chemical_4_4__DDT:matix = "SED" ;
      Chemical_4_4__DDT:units = "nanograms/gram" ;
      Chemical_4_4__DDT:_FillValue = -1. ;
      Chemical_4_4__DDT:valid_min = 0. ;
      Chemical_4_4__DDT:valid_max = 1.79769313486232e+308 ;
      Chemical_4_4__DDT:instrument = "ECDDUAL_M_Sample_dry_weight" ;
      Chemical_4_4__DDT:grid_mapping = "crs" ;
      Chemical_4_4__DDT:reference = "0074376/data/0-data/Bioeffects_Assessments/Kachemak_Bay/Data_Files/KB1_ORG.txt" ;
   double Aldrin(Sample_Site) ;
      Aldrin:long_name = "Aldrin" ;
      Aldrin:coordinates = "latitude longitude time z" ;
      Aldrin:matix = "SED" ;
      Aldrin:units = "nanograms/gram" ;
      Aldrin:_FillValue = -1. ;
      Aldrin:valid_min = 0. ;
      Aldrin:valid_max = 1.79769313486232e+308 ;
      Aldrin:instrument = "ECDDUAL_M_Sample_dry_weight" ;
      Aldrin:grid_mapping = "crs" ;
      Aldrin:reference = "0074376/data/0-data/Bioeffects_Assessments/Kachemak_Bay/Data_Files/KB1_ORG.txt" ;
   double Alpha_Chlordane(Sample_Site) ;
      Alpha_Chlordane:long_name = "Alpha-Chlordane" ;
      Alpha_Chlordane:coordinates = "latitude longitude time z" ;
      Alpha_Chlordane:matix = "SED" ;
      Alpha_Chlordane:units = "nanograms/gram" ;
      Alpha_Chlordane:_FillValue = -1. ;
      Alpha_Chlordane:valid_min = 0. ;
      Alpha_Chlordane:valid_max = 1.79769313486232e+308 ;
      Alpha_Chlordane:instrument = "ECDDUAL_M_Sample_dry_weight" ;
      Alpha_Chlordane:grid_mapping = "crs" ;
      Alpha_Chlordane:reference = "0074376/data/0-data/Bioeffects_Assessments/Kachemak_Bay/Data_Files/KB1_ORG.txt" ;
   double Alpha_Hexachlorocyclohexane(Sample_Site) ;
      Alpha_Hexachlorocyclohexane:long_name = "Alpha-Hexachlorocyclohexane" ;
      Alpha_Hexachlorocyclohexane:coordinates = "latitude longitude time z" ;
      Alpha_Hexachlorocyclohexane:matix = "SED" ;
      Alpha_Hexachlorocyclohexane:units = "nanograms/gram" ;
      Alpha_Hexachlorocyclohexane:_FillValue = -1. ;
      Alpha_Hexachlorocyclohexane:valid_min = 0. ;
      Alpha_Hexachlorocyclohexane:valid_max = 1.79769313486232e+308 ;
      Alpha_Hexachlorocyclohexane:instrument = "ECDDUAL_M_Sample_dry_weight" ;
      Alpha_Hexachlorocyclohexane:grid_mapping = "crs" ;
      Alpha_Hexachlorocyclohexane:reference = "0074376/data/0-data/Bioeffects_Assessments/Kachemak_Bay/Data_Files/KB1_ORG.txt" ;
   double Beta_Hexachlorocyclohexane(Sample_Site) ;
      Beta_Hexachlorocyclohexane:long_name = "Beta-Hexachlorocyclohexane" ;
      Beta_Hexachlorocyclohexane:coordinates = "latitude longitude time z" ;
      Beta_Hexachlorocyclohexane:matix = "SED" ;
      Beta_Hexachlorocyclohexane:units = "nanograms/gram" ;
      Beta_Hexachlorocyclohexane:_FillValue = -1. ;
      Beta_Hexachlorocyclohexane:valid_min = 0. ;
      Beta_Hexachlorocyclohexane:valid_max = 1.79769313486232e+308 ;
      Beta_Hexachlorocyclohexane:instrument = "ECDDUAL_M_Sample_dry_weight" ;
      Beta_Hexachlorocyclohexane:grid_mapping = "crs" ;
      Beta_Hexachlorocyclohexane:reference = "0074376/data/0-data/Bioeffects_Assessments/Kachemak_Bay/Data_Files/KB1_ORG.txt" ;
   double Cis_Nonachlor(Sample_Site) ;
      Cis_Nonachlor:long_name = "Cis-Nonachlor" ;
      Cis_Nonachlor:coordinates = "latitude longitude time z" ;
      Cis_Nonachlor:matix = "SED" ;
      Cis_Nonachlor:units = "nanograms/gram" ;
      Cis_Nonachlor:_FillValue = -1. ;
      Cis_Nonachlor:valid_min = 0. ;
      Cis_Nonachlor:valid_max = 1.79769313486232e+308 ;
      Cis_Nonachlor:instrument = "ECDDUAL_M_Sample_dry_weight" ;
      Cis_Nonachlor:grid_mapping = "crs" ;
      Cis_Nonachlor:reference = "0074376/data/0-data/Bioeffects_Assessments/Kachemak_Bay/Data_Files/KB1_ORG.txt" ;
   double Delta_Hexachlorocyclohexane(Sample_Site) ;
      Delta_Hexachlorocyclohexane:long_name = "Delta-Hexachlorocyclohexane" ;
      Delta_Hexachlorocyclohexane:coordinates = "latitude longitude time z" ;
      Delta_Hexachlorocyclohexane:matix = "SED" ;
      Delta_Hexachlorocyclohexane:units = "nanograms/gram" ;
      Delta_Hexachlorocyclohexane:_FillValue = -1. ;
      Delta_Hexachlorocyclohexane:valid_min = 0. ;
      Delta_Hexachlorocyclohexane:valid_max = 1.79769313486232e+308 ;
      Delta_Hexachlorocyclohexane:instrument = "ECDDUAL_M_Sample_dry_weight" ;
      Delta_Hexachlorocyclohexane:grid_mapping = "crs" ;
      Delta_Hexachlorocyclohexane:reference = "0074376/data/0-data/Bioeffects_Assessments/Kachemak_Bay/Data_Files/KB1_ORG.txt" ;
   double Dieldrin(Sample_Site) ;
      Dieldrin:long_name = "Dieldrin" ;
      Dieldrin:coordinates = "latitude longitude time z" ;
      Dieldrin:matix = "SED" ;
      Dieldrin:units = "nanograms/gram" ;
      Dieldrin:_FillValue = -1. ;
      Dieldrin:valid_min = 0. ;
      Dieldrin:valid_max = 1.79769313486232e+308 ;
      Dieldrin:instrument = "ECDDUAL_M_Sample_dry_weight" ;
      Dieldrin:grid_mapping = "crs" ;
      Dieldrin:reference = "0074376/data/0-data/Bioeffects_Assessments/Kachemak_Bay/Data_Files/KB1_ORG.txt" ;
   double Endosulfan_I(Sample_Site) ;
      Endosulfan_I:long_name = "Endosulfan I" ;
      Endosulfan_I:coordinates = "latitude longitude time z" ;
      Endosulfan_I:matix = "SED" ;
      Endosulfan_I:units = "nanograms/gram" ;
      Endosulfan_I:_FillValue = -1. ;
      Endosulfan_I:valid_min = 0. ;
      Endosulfan_I:valid_max = 1.79769313486232e+308 ;
      Endosulfan_I:instrument = "ECDDUAL_M_Sample_dry_weight" ;
      Endosulfan_I:grid_mapping = "crs" ;
      Endosulfan_I:reference = "0074376/data/0-data/Bioeffects_Assessments/Kachemak_Bay/Data_Files/KB1_ORG.txt" ;
   double Endosulfan_II(Sample_Site) ;
      Endosulfan_II:long_name = "Endosulfan II" ;
      Endosulfan_II:coordinates = "latitude longitude time z" ;
      Endosulfan_II:matix = "SED" ;
      Endosulfan_II:units = "nanograms/gram" ;
      Endosulfan_II:_FillValue = -1. ;
      Endosulfan_II:valid_min = 0. ;
      Endosulfan_II:valid_max = 1.79769313486232e+308 ;
      Endosulfan_II:instrument = "ECDDUAL_M_Sample_dry_weight" ;
      Endosulfan_II:grid_mapping = "crs" ;
      Endosulfan_II:reference = "0074376/data/0-data/Bioeffects_Assessments/Kachemak_Bay/Data_Files/KB1_ORG.txt" ;
   double Endosulfan_Sulfate(Sample_Site) ;
      Endosulfan_Sulfate:long_name = "Endosulfan Sulfate" ;
      Endosulfan_Sulfate:coordinates = "latitude longitude time z" ;
      Endosulfan_Sulfate:matix = "SED" ;
      Endosulfan_Sulfate:units = "nanograms/gram" ;
      Endosulfan_Sulfate:_FillValue = -1. ;
      Endosulfan_Sulfate:valid_min = 0. ;
      Endosulfan_Sulfate:valid_max = 1.79769313486232e+308 ;
      Endosulfan_Sulfate:instrument = "ECDDUAL_M_Sample_dry_weight" ;
      Endosulfan_Sulfate:grid_mapping = "crs" ;
      Endosulfan_Sulfate:reference = "0074376/data/0-data/Bioeffects_Assessments/Kachemak_Bay/Data_Files/KB1_ORG.txt" ;
   double Endrin(Sample_Site) ;
      Endrin:long_name = "Endrin" ;
      Endrin:coordinates = "latitude longitude time z" ;
      Endrin:matix = "SED" ;
      Endrin:units = "nanograms/gram" ;
      Endrin:_FillValue = -1. ;
      Endrin:valid_min = 0. ;
      Endrin:valid_max = 1.79769313486232e+308 ;
      Endrin:instrument = "ECDDUAL_M_Sample_dry_weight" ;
      Endrin:grid_mapping = "crs" ;
      Endrin:reference = "0074376/data/0-data/Bioeffects_Assessments/Kachemak_Bay/Data_Files/KB1_ORG.txt" ;
   double Gamma_Chlordane(Sample_Site) ;
      Gamma_Chlordane:long_name = "Gamma-Chlordane" ;
      Gamma_Chlordane:coordinates = "latitude longitude time z" ;
      Gamma_Chlordane:matix = "SED" ;
      Gamma_Chlordane:units = "nanograms/gram" ;
      Gamma_Chlordane:_FillValue = -1. ;
      Gamma_Chlordane:valid_min = 0. ;
      Gamma_Chlordane:valid_max = 1.79769313486232e+308 ;
      Gamma_Chlordane:instrument = "ECDDUAL_M_Sample_dry_weight" ;
      Gamma_Chlordane:grid_mapping = "crs" ;
      Gamma_Chlordane:reference = "0074376/data/0-data/Bioeffects_Assessments/Kachemak_Bay/Data_Files/KB1_ORG.txt" ;
   double Gamma_Hexachlorocyclohexane(Sample_Site) ;
      Gamma_Hexachlorocyclohexane:long_name = "Gamma-Hexachlorocyclohexane" ;
      Gamma_Hexachlorocyclohexane:coordinates = "latitude longitude time z" ;
      Gamma_Hexachlorocyclohexane:matix = "SED" ;
      Gamma_Hexachlorocyclohexane:units = "nanograms/gram" ;
      Gamma_Hexachlorocyclohexane:_FillValue = -1. ;
      Gamma_Hexachlorocyclohexane:valid_min = 0. ;
      Gamma_Hexachlorocyclohexane:valid_max = 1.79769313486232e+308 ;
      Gamma_Hexachlorocyclohexane:instrument = "ECDDUAL_M_Sample_dry_weight" ;
      Gamma_Hexachlorocyclohexane:grid_mapping = "crs" ;
      Gamma_Hexachlorocyclohexane:reference = "0074376/data/0-data/Bioeffects_Assessments/Kachemak_Bay/Data_Files/KB1_ORG.txt" ;
   double Heptachlor(Sample_Site) ;
      Heptachlor:long_name = "Heptachlor" ;
      Heptachlor:coordinates = "latitude longitude time z" ;
      Heptachlor:matix = "SED" ;
      Heptachlor:units = "nanograms/gram" ;
      Heptachlor:_FillValue = -1. ;
      Heptachlor:valid_min = 0. ;
      Heptachlor:valid_max = 1.79769313486232e+308 ;
      Heptachlor:instrument = "ECDDUAL_M_Sample_dry_weight" ;
      Heptachlor:grid_mapping = "crs" ;
      Heptachlor:reference = "0074376/data/0-data/Bioeffects_Assessments/Kachemak_Bay/Data_Files/KB1_ORG.txt" ;
   double Heptachlor_Epoxide(Sample_Site) ;
      Heptachlor_Epoxide:long_name = "Heptachlor-Epoxide" ;
      Heptachlor_Epoxide:coordinates = "latitude longitude time z" ;
      Heptachlor_Epoxide:matix = "SED" ;
      Heptachlor_Epoxide:units = "nanograms/gram" ;
      Heptachlor_Epoxide:_FillValue = -1. ;
      Heptachlor_Epoxide:valid_min = 0. ;
      Heptachlor_Epoxide:valid_max = 1.79769313486232e+308 ;
      Heptachlor_Epoxide:instrument = "ECDDUAL_M_Sample_dry_weight" ;
      Heptachlor_Epoxide:grid_mapping = "crs" ;
      Heptachlor_Epoxide:reference = "0074376/data/0-data/Bioeffects_Assessments/Kachemak_Bay/Data_Files/KB1_ORG.txt" ;
   double Hexachlorobenzene(Sample_Site) ;
      Hexachlorobenzene:long_name = "Hexachlorobenzene" ;
      Hexachlorobenzene:coordinates = "latitude longitude time z" ;
      Hexachlorobenzene:matix = "SED" ;
      Hexachlorobenzene:units = "nanograms/gram" ;
      Hexachlorobenzene:_FillValue = -1. ;
      Hexachlorobenzene:valid_min = 0. ;
      Hexachlorobenzene:valid_max = 1.79769313486232e+308 ;
      Hexachlorobenzene:instrument = "ECDDUAL_M_Sample_dry_weight" ;
      Hexachlorobenzene:grid_mapping = "crs" ;
      Hexachlorobenzene:reference = "0074376/data/0-data/Bioeffects_Assessments/Kachemak_Bay/Data_Files/KB1_ORG.txt" ;
   double Mirex(Sample_Site) ;
      Mirex:long_name = "Mirex" ;
      Mirex:coordinates = "latitude longitude time z" ;
      Mirex:matix = "SED" ;
      Mirex:units = "nanograms/gram" ;
      Mirex:_FillValue = -1. ;
      Mirex:valid_min = 0. ;
      Mirex:valid_max = 1.79769313486232e+308 ;
      Mirex:instrument = "ECDDUAL_M_Sample_dry_weight" ;
      Mirex:grid_mapping = "crs" ;
      Mirex:reference = "0074376/data/0-data/Bioeffects_Assessments/Kachemak_Bay/Data_Files/KB1_ORG.txt" ;
   double Oxychlordane(Sample_Site) ;
      Oxychlordane:long_name = "Oxychlordane" ;
      Oxychlordane:coordinates = "latitude longitude time z" ;
      Oxychlordane:matix = "SED" ;
      Oxychlordane:units = "nanograms/gram" ;
      Oxychlordane:_FillValue = -1. ;
      Oxychlordane:valid_min = 0. ;
      Oxychlordane:valid_max = 1.79769313486232e+308 ;
      Oxychlordane:instrument = "ECDDUAL_M_Sample_dry_weight" ;
      Oxychlordane:grid_mapping = "crs" ;
      Oxychlordane:reference = "0074376/data/0-data/Bioeffects_Assessments/Kachemak_Bay/Data_Files/KB1_ORG.txt" ;
   double PCB101_90(Sample_Site) ;
      PCB101_90:long_name = "PCB101_90" ;
      PCB101_90:coordinates = "latitude longitude time z" ;
      PCB101_90:matix = "SED" ;
      PCB101_90:units = "nanograms/gram" ;
      PCB101_90:_FillValue = -1. ;
      PCB101_90:valid_min = 0. ;
      PCB101_90:valid_max = 1.79769313486232e+308 ;
      PCB101_90:instrument = "ECDDUAL_M_Sample_dry_weight" ;
      PCB101_90:grid_mapping = "crs" ;
      PCB101_90:reference = "0074376/data/0-data/Bioeffects_Assessments/Kachemak_Bay/Data_Files/KB1_ORG.txt" ;
   double PCB105(Sample_Site) ;
      PCB105:long_name = "PCB105" ;
      PCB105:coordinates = "latitude longitude time z" ;
      PCB105:matix = "SED" ;
      PCB105:units = "nanograms/gram" ;
      PCB105:_FillValue = -1. ;
      PCB105:valid_min = 0. ;
      PCB105:valid_max = 1.79769313486232e+308 ;
      PCB105:instrument = "ECDDUAL_M_Sample_dry_weight" ;
      PCB105:grid_mapping = "crs" ;
      PCB105:reference = "0074376/data/0-data/Bioeffects_Assessments/Kachemak_Bay/Data_Files/KB1_ORG.txt" ;
   double PCB118(Sample_Site) ;
      PCB118:long_name = "PCB118" ;
      PCB118:coordinates = "latitude longitude time z" ;
      PCB118:matix = "SED" ;
      PCB118:units = "nanograms/gram" ;
      PCB118:_FillValue = -1. ;
      PCB118:valid_min = 0. ;
      PCB118:valid_max = 1.79769313486232e+308 ;
      PCB118:instrument = "ECDDUAL_M_Sample_dry_weight" ;
      PCB118:grid_mapping = "crs" ;
      PCB118:reference = "0074376/data/0-data/Bioeffects_Assessments/Kachemak_Bay/Data_Files/KB1_ORG.txt" ;
   double PCB128(Sample_Site) ;
      PCB128:long_name = "PCB128" ;
      PCB128:coordinates = "latitude longitude time z" ;
      PCB128:matix = "SED" ;
      PCB128:units = "nanograms/gram" ;
      PCB128:_FillValue = -1. ;
      PCB128:valid_min = 0. ;
      PCB128:valid_max = 1.79769313486232e+308 ;
      PCB128:instrument = "ECDDUAL_M_Sample_dry_weight" ;
      PCB128:grid_mapping = "crs" ;
      PCB128:reference = "0074376/data/0-data/Bioeffects_Assessments/Kachemak_Bay/Data_Files/KB1_ORG.txt" ;
   double PCB138_160(Sample_Site) ;
      PCB138_160:long_name = "PCB138_160" ;
      PCB138_160:coordinates = "latitude longitude time z" ;
      PCB138_160:matix = "SED" ;
      PCB138_160:units = "nanograms/gram" ;
      PCB138_160:_FillValue = -1. ;
      PCB138_160:valid_min = 0. ;
      PCB138_160:valid_max = 1.79769313486232e+308 ;
      PCB138_160:instrument = "ECDDUAL_M_Sample_dry_weight" ;
      PCB138_160:grid_mapping = "crs" ;
      PCB138_160:reference = "0074376/data/0-data/Bioeffects_Assessments/Kachemak_Bay/Data_Files/KB1_ORG.txt" ;
   double PCB146(Sample_Site) ;
      PCB146:long_name = "PCB146" ;
      PCB146:coordinates = "latitude longitude time z" ;
      PCB146:matix = "SED" ;
      PCB146:units = "nanograms/gram" ;
      PCB146:_FillValue = -1. ;
      PCB146:valid_min = 0. ;
      PCB146:valid_max = 1.79769313486232e+308 ;
      PCB146:instrument = "ECDDUAL_M_Sample_dry_weight" ;
      PCB146:grid_mapping = "crs" ;
      PCB146:reference = "0074376/data/0-data/Bioeffects_Assessments/Kachemak_Bay/Data_Files/KB1_ORG.txt" ;
   double PCB149_123(Sample_Site) ;
      PCB149_123:long_name = "PCB149_123" ;
      PCB149_123:coordinates = "latitude longitude time z" ;
      PCB149_123:matix = "SED" ;
      PCB149_123:units = "nanograms/gram" ;
      PCB149_123:_FillValue = -1. ;
      PCB149_123:valid_min = 0. ;
      PCB149_123:valid_max = 1.79769313486232e+308 ;
      PCB149_123:instrument = "ECDDUAL_M_Sample_dry_weight" ;
      PCB149_123:grid_mapping = "crs" ;
      PCB149_123:reference = "0074376/data/0-data/Bioeffects_Assessments/Kachemak_Bay/Data_Files/KB1_ORG.txt" ;
   double PCB151(Sample_Site) ;
      PCB151:long_name = "PCB151" ;
      PCB151:coordinates = "latitude longitude time z" ;
      PCB151:matix = "SED" ;
      PCB151:units = "nanograms/gram" ;
      PCB151:_FillValue = -1. ;
      PCB151:valid_min = 0. ;
      PCB151:valid_max = 1.79769313486232e+308 ;
      PCB151:instrument = "ECDDUAL_M_Sample_dry_weight" ;
      PCB151:grid_mapping = "crs" ;
      PCB151:reference = "0074376/data/0-data/Bioeffects_Assessments/Kachemak_Bay/Data_Files/KB1_ORG.txt" ;
   double PCB153_132_168(Sample_Site) ;
      PCB153_132_168:long_name = "PCB153_132_168" ;
      PCB153_132_168:coordinates = "latitude longitude time z" ;
      PCB153_132_168:matix = "SED" ;
      PCB153_132_168:units = "nanograms/gram" ;
      PCB153_132_168:_FillValue = -1. ;
      PCB153_132_168:valid_min = 0. ;
      PCB153_132_168:valid_max = 1.79769313486232e+308 ;
      PCB153_132_168:instrument = "ECDDUAL_M_Sample_dry_weight" ;
      PCB153_132_168:grid_mapping = "crs" ;
      PCB153_132_168:reference = "0074376/data/0-data/Bioeffects_Assessments/Kachemak_Bay/Data_Files/KB1_ORG.txt" ;
   double PCB156_171_202(Sample_Site) ;
      PCB156_171_202:long_name = "PCB156_171_202" ;
      PCB156_171_202:coordinates = "latitude longitude time z" ;
      PCB156_171_202:matix = "SED" ;
      PCB156_171_202:units = "nanograms/gram" ;
      PCB156_171_202:_FillValue = -1. ;
      PCB156_171_202:valid_min = 0. ;
      PCB156_171_202:valid_max = 1.79769313486232e+308 ;
      PCB156_171_202:instrument = "ECDDUAL_M_Sample_dry_weight" ;
      PCB156_171_202:grid_mapping = "crs" ;
      PCB156_171_202:reference = "0074376/data/0-data/Bioeffects_Assessments/Kachemak_Bay/Data_Files/KB1_ORG.txt" ;
   double PCB158(Sample_Site) ;
      PCB158:long_name = "PCB158" ;
      PCB158:coordinates = "latitude longitude time z" ;
      PCB158:matix = "SED" ;
      PCB158:units = "nanograms/gram" ;
      PCB158:_FillValue = -1. ;
      PCB158:valid_min = 0. ;
      PCB158:valid_max = 1.79769313486232e+308 ;
      PCB158:instrument = "ECDDUAL_M_Sample_dry_weight" ;
      PCB158:grid_mapping = "crs" ;
      PCB158:reference = "0074376/data/0-data/Bioeffects_Assessments/Kachemak_Bay/Data_Files/KB1_ORG.txt" ;
   double PCB170_190(Sample_Site) ;
      PCB170_190:long_name = "PCB170_190" ;
      PCB170_190:coordinates = "latitude longitude time z" ;
      PCB170_190:matix = "SED" ;
      PCB170_190:units = "nanograms/gram" ;
      PCB170_190:_FillValue = -1. ;
      PCB170_190:valid_min = 0. ;
      PCB170_190:valid_max = 1.79769313486232e+308 ;
      PCB170_190:instrument = "ECDDUAL_M_Sample_dry_weight" ;
      PCB170_190:grid_mapping = "crs" ;
      PCB170_190:reference = "0074376/data/0-data/Bioeffects_Assessments/Kachemak_Bay/Data_Files/KB1_ORG.txt" ;
   double PCB174(Sample_Site) ;
      PCB174:long_name = "PCB174" ;
      PCB174:coordinates = "latitude longitude time z" ;
      PCB174:matix = "SED" ;
      PCB174:units = "nanograms/gram" ;
      PCB174:_FillValue = -1. ;
      PCB174:valid_min = 0. ;
      PCB174:valid_max = 1.79769313486232e+308 ;
      PCB174:instrument = "ECDDUAL_M_Sample_dry_weight" ;
      PCB174:grid_mapping = "crs" ;
      PCB174:reference = "0074376/data/0-data/Bioeffects_Assessments/Kachemak_Bay/Data_Files/KB1_ORG.txt" ;
   double PCB18(Sample_Site) ;
      PCB18:long_name = "PCB18" ;
      PCB18:coordinates = "latitude longitude time z" ;
      PCB18:matix = "SED" ;
      PCB18:units = "nanograms/gram" ;
      PCB18:_FillValue = -1. ;
      PCB18:valid_min = 0. ;
      PCB18:valid_max = 1.79769313486232e+308 ;
      PCB18:instrument = "ECDDUAL_M_Sample_dry_weight" ;
      PCB18:grid_mapping = "crs" ;
      PCB18:reference = "0074376/data/0-data/Bioeffects_Assessments/Kachemak_Bay/Data_Files/KB1_ORG.txt" ;
   double PCB180(Sample_Site) ;
      PCB180:long_name = "PCB180" ;
      PCB180:coordinates = "latitude longitude time z" ;
      PCB180:matix = "SED" ;
      PCB180:units = "nanograms/gram" ;
      PCB180:_FillValue = -1. ;
      PCB180:valid_min = 0. ;
      PCB180:valid_max = 1.79769313486232e+308 ;
      PCB180:instrument = "ECDDUAL_M_Sample_dry_weight" ;
      PCB180:grid_mapping = "crs" ;
      PCB180:reference = "0074376/data/0-data/Bioeffects_Assessments/Kachemak_Bay/Data_Files/KB1_ORG.txt" ;
   double PCB183(Sample_Site) ;
      PCB183:long_name = "PCB183" ;
      PCB183:coordinates = "latitude longitude time z" ;
      PCB183:matix = "SED" ;
      PCB183:units = "nanograms/gram" ;
      PCB183:_FillValue = -1. ;
      PCB183:valid_min = 0. ;
      PCB183:valid_max = 1.79769313486232e+308 ;
      PCB183:instrument = "ECDDUAL_M_Sample_dry_weight" ;
      PCB183:grid_mapping = "crs" ;
      PCB183:reference = "0074376/data/0-data/Bioeffects_Assessments/Kachemak_Bay/Data_Files/KB1_ORG.txt" ;
   double PCB187(Sample_Site) ;
      PCB187:long_name = "PCB187" ;
      PCB187:coordinates = "latitude longitude time z" ;
      PCB187:matix = "SED" ;
      PCB187:units = "nanograms/gram" ;
      PCB187:_FillValue = -1. ;
      PCB187:valid_min = 0. ;
      PCB187:valid_max = 1.79769313486232e+308 ;
      PCB187:instrument = "ECDDUAL_M_Sample_dry_weight" ;
      PCB187:grid_mapping = "crs" ;
      PCB187:reference = "0074376/data/0-data/Bioeffects_Assessments/Kachemak_Bay/Data_Files/KB1_ORG.txt" ;
   double PCB194(Sample_Site) ;
      PCB194:long_name = "PCB194" ;
      PCB194:coordinates = "latitude longitude time z" ;
      PCB194:matix = "SED" ;
      PCB194:units = "nanograms/gram" ;
      PCB194:_FillValue = -1. ;
      PCB194:valid_min = 0. ;
      PCB194:valid_max = 1.79769313486232e+308 ;
      PCB194:instrument = "ECDDUAL_M_Sample_dry_weight" ;
      PCB194:grid_mapping = "crs" ;
      PCB194:reference = "0074376/data/0-data/Bioeffects_Assessments/Kachemak_Bay/Data_Files/KB1_ORG.txt" ;
   double PCB195_208(Sample_Site) ;
      PCB195_208:long_name = "PCB195_208" ;
      PCB195_208:coordinates = "latitude longitude time z" ;
      PCB195_208:matix = "SED" ;
      PCB195_208:units = "nanograms/gram" ;
      PCB195_208:_FillValue = -1. ;
      PCB195_208:valid_min = 0. ;
      PCB195_208:valid_max = 1.79769313486232e+308 ;
      PCB195_208:instrument = "ECDDUAL_M_Sample_dry_weight" ;
      PCB195_208:grid_mapping = "crs" ;
      PCB195_208:reference = "0074376/data/0-data/Bioeffects_Assessments/Kachemak_Bay/Data_Files/KB1_ORG.txt" ;
   double PCB206(Sample_Site) ;
      PCB206:long_name = "PCB206" ;
      PCB206:coordinates = "latitude longitude time z" ;
      PCB206:matix = "SED" ;
      PCB206:units = "nanograms/gram" ;
      PCB206:_FillValue = -1. ;
      PCB206:valid_min = 0. ;
      PCB206:valid_max = 1.79769313486232e+308 ;
      PCB206:instrument = "ECDDUAL_M_Sample_dry_weight" ;
      PCB206:grid_mapping = "crs" ;
      PCB206:reference = "0074376/data/0-data/Bioeffects_Assessments/Kachemak_Bay/Data_Files/KB1_ORG.txt" ;
   double PCB209(Sample_Site) ;
      PCB209:long_name = "PCB209" ;
      PCB209:coordinates = "latitude longitude time z" ;
      PCB209:matix = "SED" ;
      PCB209:units = "nanograms/gram" ;
      PCB209:_FillValue = -1. ;
      PCB209:valid_min = 0. ;
      PCB209:valid_max = 1.79769313486232e+308 ;
      PCB209:instrument = "ECDDUAL_M_Sample_dry_weight" ;
      PCB209:grid_mapping = "crs" ;
      PCB209:reference = "0074376/data/0-data/Bioeffects_Assessments/Kachemak_Bay/Data_Files/KB1_ORG.txt" ;
   double PCB28(Sample_Site) ;
      PCB28:long_name = "PCB28" ;
      PCB28:coordinates = "latitude longitude time z" ;
      PCB28:matix = "SED" ;
      PCB28:units = "nanograms/gram" ;
      PCB28:_FillValue = -1. ;
      PCB28:valid_min = 0. ;
      PCB28:valid_max = 1.79769313486232e+308 ;
      PCB28:instrument = "ECDDUAL_M_Sample_dry_weight" ;
      PCB28:grid_mapping = "crs" ;
      PCB28:reference = "0074376/data/0-data/Bioeffects_Assessments/Kachemak_Bay/Data_Files/KB1_ORG.txt" ;
   double PCB29(Sample_Site) ;
      PCB29:long_name = "PCB29" ;
      PCB29:coordinates = "latitude longitude time z" ;
      PCB29:matix = "SED" ;
      PCB29:units = "nanograms/gram" ;
      PCB29:_FillValue = -1. ;
      PCB29:valid_min = 0. ;
      PCB29:valid_max = 1.79769313486232e+308 ;
      PCB29:instrument = "ECDDUAL_M_Sample_dry_weight" ;
      PCB29:grid_mapping = "crs" ;
      PCB29:reference = "0074376/data/0-data/Bioeffects_Assessments/Kachemak_Bay/Data_Files/KB1_ORG.txt" ;
   double PCB31(Sample_Site) ;
      PCB31:long_name = "PCB31" ;
      PCB31:coordinates = "latitude longitude time z" ;
      PCB31:matix = "SED" ;
      PCB31:units = "nanograms/gram" ;
      PCB31:_FillValue = -1. ;
      PCB31:valid_min = 0. ;
      PCB31:valid_max = 1.79769313486232e+308 ;
      PCB31:instrument = "ECDDUAL_M_Sample_dry_weight" ;
      PCB31:grid_mapping = "crs" ;
      PCB31:reference = "0074376/data/0-data/Bioeffects_Assessments/Kachemak_Bay/Data_Files/KB1_ORG.txt" ;
   double PCB44(Sample_Site) ;
      PCB44:long_name = "PCB44" ;
      PCB44:coordinates = "latitude longitude time z" ;
      PCB44:matix = "SED" ;
      PCB44:units = "nanograms/gram" ;
      PCB44:_FillValue = -1. ;
      PCB44:valid_min = 0. ;
      PCB44:valid_max = 1.79769313486232e+308 ;
      PCB44:instrument = "ECDDUAL_M_Sample_dry_weight" ;
      PCB44:grid_mapping = "crs" ;
      PCB44:reference = "0074376/data/0-data/Bioeffects_Assessments/Kachemak_Bay/Data_Files/KB1_ORG.txt" ;
   double PCB45(Sample_Site) ;
      PCB45:long_name = "PCB45" ;
      PCB45:coordinates = "latitude longitude time z" ;
      PCB45:matix = "SED" ;
      PCB45:units = "nanograms/gram" ;
      PCB45:_FillValue = -1. ;
      PCB45:valid_min = 0. ;
      PCB45:valid_max = 1.79769313486232e+308 ;
      PCB45:instrument = "ECDDUAL_M_Sample_dry_weight" ;
      PCB45:grid_mapping = "crs" ;
      PCB45:reference = "0074376/data/0-data/Bioeffects_Assessments/Kachemak_Bay/Data_Files/KB1_ORG.txt" ;
   double PCB49(Sample_Site) ;
      PCB49:long_name = "PCB49" ;
      PCB49:coordinates = "latitude longitude time z" ;
      PCB49:matix = "SED" ;
      PCB49:units = "nanograms/gram" ;
      PCB49:_FillValue = -1. ;
      PCB49:valid_min = 0. ;
      PCB49:valid_max = 1.79769313486232e+308 ;
      PCB49:instrument = "ECDDUAL_M_Sample_dry_weight" ;
      PCB49:grid_mapping = "crs" ;
      PCB49:reference = "0074376/data/0-data/Bioeffects_Assessments/Kachemak_Bay/Data_Files/KB1_ORG.txt" ;
   double PCB52(Sample_Site) ;
      PCB52:long_name = "PCB52" ;
      PCB52:coordinates = "latitude longitude time z" ;
      PCB52:matix = "SED" ;
      PCB52:units = "nanograms/gram" ;
      PCB52:_FillValue = -1. ;
      PCB52:valid_min = 0. ;
      PCB52:valid_max = 1.79769313486232e+308 ;
      PCB52:instrument = "ECDDUAL_M_Sample_dry_weight" ;
      PCB52:grid_mapping = "crs" ;
      PCB52:reference = "0074376/data/0-data/Bioeffects_Assessments/Kachemak_Bay/Data_Files/KB1_ORG.txt" ;
   double PCB56_60(Sample_Site) ;
      PCB56_60:long_name = "PCB56_60" ;
      PCB56_60:coordinates = "latitude longitude time z" ;
      PCB56_60:matix = "SED" ;
      PCB56_60:units = "nanograms/gram" ;
      PCB56_60:_FillValue = -1. ;
      PCB56_60:valid_min = 0. ;
      PCB56_60:valid_max = 1.79769313486232e+308 ;
      PCB56_60:instrument = "ECDDUAL_M_Sample_dry_weight" ;
      PCB56_60:grid_mapping = "crs" ;
      PCB56_60:reference = "0074376/data/0-data/Bioeffects_Assessments/Kachemak_Bay/Data_Files/KB1_ORG.txt" ;
   double PCB66(Sample_Site) ;
      PCB66:long_name = "PCB66" ;
      PCB66:coordinates = "latitude longitude time z" ;
      PCB66:matix = "SED" ;
      PCB66:units = "nanograms/gram" ;
      PCB66:_FillValue = -1. ;
      PCB66:valid_min = 0. ;
      PCB66:valid_max = 1.79769313486232e+308 ;
      PCB66:instrument = "ECDDUAL_M_Sample_dry_weight" ;
      PCB66:grid_mapping = "crs" ;
      PCB66:reference = "0074376/data/0-data/Bioeffects_Assessments/Kachemak_Bay/Data_Files/KB1_ORG.txt" ;
   double PCB70(Sample_Site) ;
      PCB70:long_name = "PCB70" ;
      PCB70:coordinates = "latitude longitude time z" ;
      PCB70:matix = "SED" ;
      PCB70:units = "nanograms/gram" ;
      PCB70:_FillValue = -1. ;
      PCB70:valid_min = 0. ;
      PCB70:valid_max = 1.79769313486232e+308 ;
      PCB70:instrument = "ECDDUAL_M_Sample_dry_weight" ;
      PCB70:grid_mapping = "crs" ;
      PCB70:reference = "0074376/data/0-data/Bioeffects_Assessments/Kachemak_Bay/Data_Files/KB1_ORG.txt" ;
   double PCB74_61(Sample_Site) ;
      PCB74_61:long_name = "PCB74_61" ;
      PCB74_61:coordinates = "latitude longitude time z" ;
      PCB74_61:matix = "SED" ;
      PCB74_61:units = "nanograms/gram" ;
      PCB74_61:_FillValue = -1. ;
      PCB74_61:valid_min = 0. ;
      PCB74_61:valid_max = 1.79769313486232e+308 ;
      PCB74_61:instrument = "ECDDUAL_M_Sample_dry_weight" ;
      PCB74_61:grid_mapping = "crs" ;
      PCB74_61:reference = "0074376/data/0-data/Bioeffects_Assessments/Kachemak_Bay/Data_Files/KB1_ORG.txt" ;
   double PCB87_115(Sample_Site) ;
      PCB87_115:long_name = "PCB87_115" ;
      PCB87_115:coordinates = "latitude longitude time z" ;
      PCB87_115:matix = "SED" ;
      PCB87_115:units = "nanograms/gram" ;
      PCB87_115:_FillValue = -1. ;
      PCB87_115:valid_min = 0. ;
      PCB87_115:valid_max = 1.79769313486232e+308 ;
      PCB87_115:instrument = "ECDDUAL_M_Sample_dry_weight" ;
      PCB87_115:grid_mapping = "crs" ;
      PCB87_115:reference = "0074376/data/0-data/Bioeffects_Assessments/Kachemak_Bay/Data_Files/KB1_ORG.txt" ;
   double PCB8_5(Sample_Site) ;
      PCB8_5:long_name = "PCB8_5" ;
      PCB8_5:coordinates = "latitude longitude time z" ;
      PCB8_5:matix = "SED" ;
      PCB8_5:units = "nanograms/gram" ;
      PCB8_5:_FillValue = -1. ;
      PCB8_5:valid_min = 0. ;
      PCB8_5:valid_max = 1.79769313486232e+308 ;
      PCB8_5:instrument = "ECDDUAL_M_Sample_dry_weight" ;
      PCB8_5:grid_mapping = "crs" ;
      PCB8_5:reference = "0074376/data/0-data/Bioeffects_Assessments/Kachemak_Bay/Data_Files/KB1_ORG.txt" ;
   double PCB95(Sample_Site) ;
      PCB95:long_name = "PCB95" ;
      PCB95:coordinates = "latitude longitude time z" ;
      PCB95:matix = "SED" ;
      PCB95:units = "nanograms/gram" ;
      PCB95:_FillValue = -1. ;
      PCB95:valid_min = 0. ;
      PCB95:valid_max = 1.79769313486232e+308 ;
      PCB95:instrument = "ECDDUAL_M_Sample_dry_weight" ;
      PCB95:grid_mapping = "crs" ;
      PCB95:reference = "0074376/data/0-data/Bioeffects_Assessments/Kachemak_Bay/Data_Files/KB1_ORG.txt" ;
   double PCB99(Sample_Site) ;
      PCB99:long_name = "PCB99" ;
      PCB99:coordinates = "latitude longitude time z" ;
      PCB99:matix = "SED" ;
      PCB99:units = "nanograms/gram" ;
      PCB99:_FillValue = -1. ;
      PCB99:valid_min = 0. ;
      PCB99:valid_max = 1.79769313486232e+308 ;
      PCB99:instrument = "ECDDUAL_M_Sample_dry_weight" ;
      PCB99:grid_mapping = "crs" ;
      PCB99:reference = "0074376/data/0-data/Bioeffects_Assessments/Kachemak_Bay/Data_Files/KB1_ORG.txt" ;
   double Pentachloroanisole(Sample_Site) ;
      Pentachloroanisole:long_name = "Pentachloroanisole" ;
      Pentachloroanisole:coordinates = "latitude longitude time z" ;
      Pentachloroanisole:matix = "SED" ;
      Pentachloroanisole:units = "nanograms/gram" ;
      Pentachloroanisole:_FillValue = -1. ;
      Pentachloroanisole:valid_min = 0. ;
      Pentachloroanisole:valid_max = 1.79769313486232e+308 ;
      Pentachloroanisole:instrument = "ECDDUAL_M_Sample_dry_weight" ;
      Pentachloroanisole:grid_mapping = "crs" ;
      Pentachloroanisole:reference = "0074376/data/0-data/Bioeffects_Assessments/Kachemak_Bay/Data_Files/KB1_ORG.txt" ;
   double Pentachlorobenzene(Sample_Site) ;
      Pentachlorobenzene:long_name = "Pentachlorobenzene" ;
      Pentachlorobenzene:coordinates = "latitude longitude time z" ;
      Pentachlorobenzene:matix = "SED" ;
      Pentachlorobenzene:units = "nanograms/gram" ;
      Pentachlorobenzene:_FillValue = -1. ;
      Pentachlorobenzene:valid_min = 0. ;
      Pentachlorobenzene:valid_max = 1.79769313486232e+308 ;
      Pentachlorobenzene:instrument = "ECDDUAL_M_Sample_dry_weight" ;
      Pentachlorobenzene:grid_mapping = "crs" ;
      Pentachlorobenzene:reference = "0074376/data/0-data/Bioeffects_Assessments/Kachemak_Bay/Data_Files/KB1_ORG.txt" ;
   double ECDDUAL_M_Sample_dry_weight(Sample_Site) ;
      ECDDUAL_M_Sample_dry_weight:long_name = "Sample dry weight" ;
      ECDDUAL_M_Sample_dry_weight:coordinates = "latitude longitude time z" ;
      ECDDUAL_M_Sample_dry_weight:matix = "SED" ;
      ECDDUAL_M_Sample_dry_weight:units = "gram" ;
      ECDDUAL_M_Sample_dry_weight:_FillValue = -1. ;
      ECDDUAL_M_Sample_dry_weight:valid_min = 0. ;
      ECDDUAL_M_Sample_dry_weight:valid_max = 1.79769313486232e+308 ;
      ECDDUAL_M_Sample_dry_weight:instrument = "ECDDUAL_M" ;
      ECDDUAL_M_Sample_dry_weight:grid_mapping = "crs" ;
      ECDDUAL_M_Sample_dry_weight:reference = "0074376/data/0-data/Bioeffects_Assessments/Kachemak_Bay/Data_Files/KB1_ORG.txt" ;
   double ECDDUAL_M_Sample_percent_dry_weight(Sample_Site) ;
      ECDDUAL_M_Sample_percent_dry_weight:long_name = "Sample percent dry weight" ;
      ECDDUAL_M_Sample_percent_dry_weight:coordinates = "latitude longitude time z" ;
      ECDDUAL_M_Sample_percent_dry_weight:matix = "SED" ;
      ECDDUAL_M_Sample_percent_dry_weight:units = "percent" ;
      ECDDUAL_M_Sample_percent_dry_weight:_FillValue = -1. ;
      ECDDUAL_M_Sample_percent_dry_weight:valid_min = 0. ;
      ECDDUAL_M_Sample_percent_dry_weight:valid_max = 100. ;
      ECDDUAL_M_Sample_percent_dry_weight:instrument = "ECDDUAL_M" ;
      ECDDUAL_M_Sample_percent_dry_weight:grid_mapping = "crs" ;
      ECDDUAL_M_Sample_percent_dry_weight:reference = "0074376/data/0-data/Bioeffects_Assessments/Kachemak_Bay/Data_Files/KB1_ORG.txt" ;
   double ECDDUAL_M_Sample_percent_wet_weight(Sample_Site) ;
      ECDDUAL_M_Sample_percent_wet_weight:long_name = "Sample percent wet weight" ;
      ECDDUAL_M_Sample_percent_wet_weight:coordinates = "latitude longitude time z" ;
      ECDDUAL_M_Sample_percent_wet_weight:matix = "SED" ;
      ECDDUAL_M_Sample_percent_wet_weight:units = "percent" ;
      ECDDUAL_M_Sample_percent_wet_weight:_FillValue = -1. ;
      ECDDUAL_M_Sample_percent_wet_weight:valid_min = 0. ;
      ECDDUAL_M_Sample_percent_wet_weight:valid_max = 100. ;
      ECDDUAL_M_Sample_percent_wet_weight:instrument = "ECDDUAL_M" ;
      ECDDUAL_M_Sample_percent_wet_weight:grid_mapping = "crs" ;
      ECDDUAL_M_Sample_percent_wet_weight:reference = "0074376/data/0-data/Bioeffects_Assessments/Kachemak_Bay/Data_Files/KB1_ORG.txt" ;
   double ECDDUAL_M_Sample_wet_weight(Sample_Site) ;
      ECDDUAL_M_Sample_wet_weight:long_name = "Sample wet weight" ;
      ECDDUAL_M_Sample_wet_weight:coordinates = "latitude longitude time z" ;
      ECDDUAL_M_Sample_wet_weight:matix = "SED" ;
      ECDDUAL_M_Sample_wet_weight:units = "gram" ;
      ECDDUAL_M_Sample_wet_weight:_FillValue = -1. ;
      ECDDUAL_M_Sample_wet_weight:valid_min = 0. ;
      ECDDUAL_M_Sample_wet_weight:valid_max = 1.79769313486232e+308 ;
      ECDDUAL_M_Sample_wet_weight:instrument = "ECDDUAL_M" ;
      ECDDUAL_M_Sample_wet_weight:grid_mapping = "crs" ;
      ECDDUAL_M_Sample_wet_weight:reference = "0074376/data/0-data/Bioeffects_Assessments/Kachemak_Bay/Data_Files/KB1_ORG.txt" ;
   double Trans_Nonachlor(Sample_Site) ;
      Trans_Nonachlor:long_name = "Trans-Nonachlor" ;
      Trans_Nonachlor:coordinates = "latitude longitude time z" ;
      Trans_Nonachlor:matix = "SED" ;
      Trans_Nonachlor:units = "nanograms/gram" ;
      Trans_Nonachlor:_FillValue = -1. ;
      Trans_Nonachlor:valid_min = 0. ;
      Trans_Nonachlor:valid_max = 1.79769313486232e+308 ;
      Trans_Nonachlor:instrument = "ECDDUAL_M_Sample_dry_weight" ;
      Trans_Nonachlor:grid_mapping = "crs" ;
      Trans_Nonachlor:reference = "0074376/data/0-data/Bioeffects_Assessments/Kachemak_Bay/Data_Files/KB1_ORG.txt" ;
   double Clay___Chemistry_Sample(Sample_Site) ;
      Clay___Chemistry_Sample:long_name = "Clay - Chemistry Sample" ;
      Clay___Chemistry_Sample:coordinates = "latitude longitude time z" ;
      Clay___Chemistry_Sample:matix = "SED" ;
      Clay___Chemistry_Sample:units = "percent" ;
      Clay___Chemistry_Sample:_FillValue = -1. ;
      Clay___Chemistry_Sample:valid_min = 0. ;
      Clay___Chemistry_Sample:valid_max = 100. ;
      Clay___Chemistry_Sample:instrument = "GS" ;
      Clay___Chemistry_Sample:grid_mapping = "crs" ;
      Clay___Chemistry_Sample:reference = "0074376/data/0-data/Bioeffects_Assessments/Kachemak_Bay/Data_Files/KB1_ORG.txt" ;
   double Gravel___Chemistry_Sample(Sample_Site) ;
      Gravel___Chemistry_Sample:long_name = "Gravel - Chemistry Sample" ;
      Gravel___Chemistry_Sample:coordinates = "latitude longitude time z" ;
      Gravel___Chemistry_Sample:matix = "SED" ;
      Gravel___Chemistry_Sample:units = "percent" ;
      Gravel___Chemistry_Sample:_FillValue = -1. ;
      Gravel___Chemistry_Sample:valid_min = 0. ;
      Gravel___Chemistry_Sample:valid_max = 100. ;
      Gravel___Chemistry_Sample:instrument = "GS" ;
      Gravel___Chemistry_Sample:grid_mapping = "crs" ;
      Gravel___Chemistry_Sample:reference = "0074376/data/0-data/Bioeffects_Assessments/Kachemak_Bay/Data_Files/KB1_ORG.txt" ;
   double GS_Sample_dry_weight(Sample_Site) ;
      GS_Sample_dry_weight:long_name = "Sample dry weight" ;
      GS_Sample_dry_weight:coordinates = "latitude longitude time z" ;
      GS_Sample_dry_weight:matix = "SED" ;
      GS_Sample_dry_weight:units = "gram" ;
      GS_Sample_dry_weight:_FillValue = -1. ;
      GS_Sample_dry_weight:valid_min = 0. ;
      GS_Sample_dry_weight:valid_max = 1.79769313486232e+308 ;
      GS_Sample_dry_weight:instrument = "GS" ;
      GS_Sample_dry_weight:grid_mapping = "crs" ;
      GS_Sample_dry_weight:reference = "0074376/data/0-data/Bioeffects_Assessments/Kachemak_Bay/Data_Files/KB1_ORG.txt" ;
   double Sand___Chemistry_Sample(Sample_Site) ;
      Sand___Chemistry_Sample:long_name = "Sand - Chemistry Sample" ;
      Sand___Chemistry_Sample:coordinates = "latitude longitude time z" ;
      Sand___Chemistry_Sample:matix = "SED" ;
      Sand___Chemistry_Sample:units = "percent" ;
      Sand___Chemistry_Sample:_FillValue = -1. ;
      Sand___Chemistry_Sample:valid_min = 0. ;
      Sand___Chemistry_Sample:valid_max = 100. ;
      Sand___Chemistry_Sample:instrument = "GS" ;
      Sand___Chemistry_Sample:grid_mapping = "crs" ;
      Sand___Chemistry_Sample:reference = "0074376/data/0-data/Bioeffects_Assessments/Kachemak_Bay/Data_Files/KB1_ORG.txt" ;
   double Silt___Chemistry_Sample(Sample_Site) ;
      Silt___Chemistry_Sample:long_name = "Silt - Chemistry Sample" ;
      Silt___Chemistry_Sample:coordinates = "latitude longitude time z" ;
      Silt___Chemistry_Sample:matix = "SED" ;
      Silt___Chemistry_Sample:units = "percent" ;
      Silt___Chemistry_Sample:_FillValue = -1. ;
      Silt___Chemistry_Sample:valid_min = 0. ;
      Silt___Chemistry_Sample:valid_max = 100. ;
      Silt___Chemistry_Sample:instrument = "GS" ;
      Silt___Chemistry_Sample:grid_mapping = "crs" ;
      Silt___Chemistry_Sample:reference = "0074376/data/0-data/Bioeffects_Assessments/Kachemak_Bay/Data_Files/KB1_ORG.txt" ;
   double Hexylation_Sample_dry_weight(Sample_Site) ;
      Hexylation_Sample_dry_weight:long_name = "Sample dry weight" ;
      Hexylation_Sample_dry_weight:coordinates = "latitude longitude time z" ;
      Hexylation_Sample_dry_weight:matix = "SED" ;
      Hexylation_Sample_dry_weight:units = "gram" ;
      Hexylation_Sample_dry_weight:_FillValue = -1. ;
      Hexylation_Sample_dry_weight:valid_min = 0. ;
      Hexylation_Sample_dry_weight:valid_max = 1.79769313486232e+308 ;
      Hexylation_Sample_dry_weight:instrument = "Hexylation" ;
      Hexylation_Sample_dry_weight:grid_mapping = "crs" ;
      Hexylation_Sample_dry_weight:reference = "0074376/data/0-data/Bioeffects_Assessments/Kachemak_Bay/Data_Files/KB1_ORG.txt" ;
   double Hexylation_Sample_percent_dry_weight(Sample_Site) ;
      Hexylation_Sample_percent_dry_weight:long_name = "Sample percent dry weight" ;
      Hexylation_Sample_percent_dry_weight:coordinates = "latitude longitude time z" ;
      Hexylation_Sample_percent_dry_weight:matix = "SED" ;
      Hexylation_Sample_percent_dry_weight:units = "percent" ;
      Hexylation_Sample_percent_dry_weight:_FillValue = -1. ;
      Hexylation_Sample_percent_dry_weight:valid_min = 0. ;
      Hexylation_Sample_percent_dry_weight:valid_max = 100. ;
      Hexylation_Sample_percent_dry_weight:instrument = "Hexylation" ;
      Hexylation_Sample_percent_dry_weight:grid_mapping = "crs" ;
      Hexylation_Sample_percent_dry_weight:reference = "0074376/data/0-data/Bioeffects_Assessments/Kachemak_Bay/Data_Files/KB1_ORG.txt" ;
   double Hexylation_Sample_percent_wet_weight(Sample_Site) ;
      Hexylation_Sample_percent_wet_weight:long_name = "Sample percent wet weight" ;
      Hexylation_Sample_percent_wet_weight:coordinates = "latitude longitude time z" ;
      Hexylation_Sample_percent_wet_weight:matix = "SED" ;
      Hexylation_Sample_percent_wet_weight:units = "percent" ;
      Hexylation_Sample_percent_wet_weight:_FillValue = -1. ;
      Hexylation_Sample_percent_wet_weight:valid_min = 0. ;
      Hexylation_Sample_percent_wet_weight:valid_max = 100. ;
      Hexylation_Sample_percent_wet_weight:instrument = "Hexylation" ;
      Hexylation_Sample_percent_wet_weight:grid_mapping = "crs" ;
      Hexylation_Sample_percent_wet_weight:reference = "0074376/data/0-data/Bioeffects_Assessments/Kachemak_Bay/Data_Files/KB1_ORG.txt" ;
   double Hexylation_Sample_wet_weight(Sample_Site) ;
      Hexylation_Sample_wet_weight:long_name = "Sample wet weight" ;
      Hexylation_Sample_wet_weight:coordinates = "latitude longitude time z" ;
      Hexylation_Sample_wet_weight:matix = "SED" ;
      Hexylation_Sample_wet_weight:units = "gram" ;
      Hexylation_Sample_wet_weight:_FillValue = -1. ;
      Hexylation_Sample_wet_weight:valid_min = 0. ;
      Hexylation_Sample_wet_weight:valid_max = 1.79769313486232e+308 ;
      Hexylation_Sample_wet_weight:instrument = "Hexylation" ;
      Hexylation_Sample_wet_weight:grid_mapping = "crs" ;
      Hexylation_Sample_wet_weight:reference = "0074376/data/0-data/Bioeffects_Assessments/Kachemak_Bay/Data_Files/KB1_ORG.txt" ;
   double Tributyltin(Sample_Site) ;
      Tributyltin:long_name = "Tributyltin" ;
      Tributyltin:coordinates = "latitude longitude time z" ;
      Tributyltin:matix = "SED" ;
      Tributyltin:units = "ngram/gram" ;
      Tributyltin:_FillValue = -1. ;
      Tributyltin:valid_min = 0. ;
      Tributyltin:valid_max = 1.79769313486232e+308 ;
      Tributyltin:instrument = "Hexylation_Sample_dry_weight" ;
      Tributyltin:grid_mapping = "crs" ;
      Tributyltin:reference = "0074376/data/0-data/Bioeffects_Assessments/Kachemak_Bay/Data_Files/KB1_ORG.txt" ;
   double Chemical_1_6_7_Trimethylnaphthalene(Sample_Site) ;
      Chemical_1_6_7_Trimethylnaphthalene:long_name = "1,6,7-Trimethylnaphthalene" ;
      Chemical_1_6_7_Trimethylnaphthalene:coordinates = "latitude longitude time z" ;
      Chemical_1_6_7_Trimethylnaphthalene:matix = "SED" ;
      Chemical_1_6_7_Trimethylnaphthalene:units = "nanograms/gram" ;
      Chemical_1_6_7_Trimethylnaphthalene:_FillValue = -1. ;
      Chemical_1_6_7_Trimethylnaphthalene:valid_min = 0. ;
      Chemical_1_6_7_Trimethylnaphthalene:valid_max = 1.79769313486232e+308 ;
      Chemical_1_6_7_Trimethylnaphthalene:instrument = "PAH_2002_Sample_dry_weight" ;
      Chemical_1_6_7_Trimethylnaphthalene:grid_mapping = "crs" ;
      Chemical_1_6_7_Trimethylnaphthalene:reference = "0074376/data/0-data/Bioeffects_Assessments/Kachemak_Bay/Data_Files/KB1_ORG.txt" ;
   double Chemical_1_Methylnaphthalene(Sample_Site) ;
      Chemical_1_Methylnaphthalene:long_name = "1-Methylnaphthalene" ;
      Chemical_1_Methylnaphthalene:coordinates = "latitude longitude time z" ;
      Chemical_1_Methylnaphthalene:matix = "SED" ;
      Chemical_1_Methylnaphthalene:units = "nanograms/gram" ;
      Chemical_1_Methylnaphthalene:_FillValue = -1. ;
      Chemical_1_Methylnaphthalene:valid_min = 0. ;
      Chemical_1_Methylnaphthalene:valid_max = 1.79769313486232e+308 ;
      Chemical_1_Methylnaphthalene:instrument = "PAH_2002_Sample_dry_weight" ;
      Chemical_1_Methylnaphthalene:grid_mapping = "crs" ;
      Chemical_1_Methylnaphthalene:reference = "0074376/data/0-data/Bioeffects_Assessments/Kachemak_Bay/Data_Files/KB1_ORG.txt" ;
   double Chemical_1_Methylphenanthrene(Sample_Site) ;
      Chemical_1_Methylphenanthrene:long_name = "1-Methylphenanthrene" ;
      Chemical_1_Methylphenanthrene:coordinates = "latitude longitude time z" ;
      Chemical_1_Methylphenanthrene:matix = "SED" ;
      Chemical_1_Methylphenanthrene:units = "nanograms/gram" ;
      Chemical_1_Methylphenanthrene:_FillValue = -1. ;
      Chemical_1_Methylphenanthrene:valid_min = 0. ;
      Chemical_1_Methylphenanthrene:valid_max = 1.79769313486232e+308 ;
      Chemical_1_Methylphenanthrene:instrument = "PAH_2002_Sample_dry_weight" ;
      Chemical_1_Methylphenanthrene:grid_mapping = "crs" ;
      Chemical_1_Methylphenanthrene:reference = "0074376/data/0-data/Bioeffects_Assessments/Kachemak_Bay/Data_Files/KB1_ORG.txt" ;
   double Chemical_2_6_Dimethylnaphthalene(Sample_Site) ;
      Chemical_2_6_Dimethylnaphthalene:long_name = "2,6-Dimethylnaphthalene" ;
      Chemical_2_6_Dimethylnaphthalene:coordinates = "latitude longitude time z" ;
      Chemical_2_6_Dimethylnaphthalene:matix = "SED" ;
      Chemical_2_6_Dimethylnaphthalene:units = "nanograms/gram" ;
      Chemical_2_6_Dimethylnaphthalene:_FillValue = -1. ;
      Chemical_2_6_Dimethylnaphthalene:valid_min = 0. ;
      Chemical_2_6_Dimethylnaphthalene:valid_max = 1.79769313486232e+308 ;
      Chemical_2_6_Dimethylnaphthalene:instrument = "PAH_2002_Sample_dry_weight" ;
      Chemical_2_6_Dimethylnaphthalene:grid_mapping = "crs" ;
      Chemical_2_6_Dimethylnaphthalene:reference = "0074376/data/0-data/Bioeffects_Assessments/Kachemak_Bay/Data_Files/KB1_ORG.txt" ;
   double Chemical_2_Methylnaphthalene(Sample_Site) ;
      Chemical_2_Methylnaphthalene:long_name = "2-Methylnaphthalene" ;
      Chemical_2_Methylnaphthalene:coordinates = "latitude longitude time z" ;
      Chemical_2_Methylnaphthalene:matix = "SED" ;
      Chemical_2_Methylnaphthalene:units = "nanograms/gram" ;
      Chemical_2_Methylnaphthalene:_FillValue = -1. ;
      Chemical_2_Methylnaphthalene:valid_min = 0. ;
      Chemical_2_Methylnaphthalene:valid_max = 1.79769313486232e+308 ;
      Chemical_2_Methylnaphthalene:instrument = "PAH_2002_Sample_dry_weight" ;
      Chemical_2_Methylnaphthalene:grid_mapping = "crs" ;
      Chemical_2_Methylnaphthalene:reference = "0074376/data/0-data/Bioeffects_Assessments/Kachemak_Bay/Data_Files/KB1_ORG.txt" ;
   double Acenaphthene(Sample_Site) ;
      Acenaphthene:long_name = "Acenaphthene" ;
      Acenaphthene:coordinates = "latitude longitude time z" ;
      Acenaphthene:matix = "SED" ;
      Acenaphthene:units = "nanograms/gram" ;
      Acenaphthene:_FillValue = -1. ;
      Acenaphthene:valid_min = 0. ;
      Acenaphthene:valid_max = 1.79769313486232e+308 ;
      Acenaphthene:instrument = "PAH_2002_Sample_dry_weight" ;
      Acenaphthene:grid_mapping = "crs" ;
      Acenaphthene:reference = "0074376/data/0-data/Bioeffects_Assessments/Kachemak_Bay/Data_Files/KB1_ORG.txt" ;
   double Acenaphthylene(Sample_Site) ;
      Acenaphthylene:long_name = "Acenaphthylene" ;
      Acenaphthylene:coordinates = "latitude longitude time z" ;
      Acenaphthylene:matix = "SED" ;
      Acenaphthylene:units = "nanograms/gram" ;
      Acenaphthylene:_FillValue = -1. ;
      Acenaphthylene:valid_min = 0. ;
      Acenaphthylene:valid_max = 1.79769313486232e+308 ;
      Acenaphthylene:instrument = "PAH_2002_Sample_dry_weight" ;
      Acenaphthylene:grid_mapping = "crs" ;
      Acenaphthylene:reference = "0074376/data/0-data/Bioeffects_Assessments/Kachemak_Bay/Data_Files/KB1_ORG.txt" ;
   double Anthracene(Sample_Site) ;
      Anthracene:long_name = "Anthracene" ;
      Anthracene:coordinates = "latitude longitude time z" ;
      Anthracene:matix = "SED" ;
      Anthracene:units = "nanograms/gram" ;
      Anthracene:_FillValue = -1. ;
      Anthracene:valid_min = 0. ;
      Anthracene:valid_max = 1.79769313486232e+308 ;
      Anthracene:instrument = "PAH_2002_Sample_dry_weight" ;
      Anthracene:grid_mapping = "crs" ;
      Anthracene:reference = "0074376/data/0-data/Bioeffects_Assessments/Kachemak_Bay/Data_Files/KB1_ORG.txt" ;
   double Benz_a_anthracene(Sample_Site) ;
      Benz_a_anthracene:long_name = "Benz[a]anthracene" ;
      Benz_a_anthracene:coordinates = "latitude longitude time z" ;
      Benz_a_anthracene:matix = "SED" ;
      Benz_a_anthracene:units = "nanograms/gram" ;
      Benz_a_anthracene:_FillValue = -1. ;
      Benz_a_anthracene:valid_min = 0. ;
      Benz_a_anthracene:valid_max = 1.79769313486232e+308 ;
      Benz_a_anthracene:instrument = "PAH_2002_Sample_dry_weight" ;
      Benz_a_anthracene:grid_mapping = "crs" ;
      Benz_a_anthracene:reference = "0074376/data/0-data/Bioeffects_Assessments/Kachemak_Bay/Data_Files/KB1_ORG.txt" ;
   double Benzo_a_pyrene(Sample_Site) ;
      Benzo_a_pyrene:long_name = "Benzo[a]pyrene" ;
      Benzo_a_pyrene:coordinates = "latitude longitude time z" ;
      Benzo_a_pyrene:matix = "SED" ;
      Benzo_a_pyrene:units = "nanograms/gram" ;
      Benzo_a_pyrene:_FillValue = -1. ;
      Benzo_a_pyrene:valid_min = 0. ;
      Benzo_a_pyrene:valid_max = 1.79769313486232e+308 ;
      Benzo_a_pyrene:instrument = "PAH_2002_Sample_dry_weight" ;
      Benzo_a_pyrene:grid_mapping = "crs" ;
      Benzo_a_pyrene:reference = "0074376/data/0-data/Bioeffects_Assessments/Kachemak_Bay/Data_Files/KB1_ORG.txt" ;
   double Benzo_b_fluoranthene(Sample_Site) ;
      Benzo_b_fluoranthene:long_name = "Benzo[b]fluoranthene" ;
      Benzo_b_fluoranthene:coordinates = "latitude longitude time z" ;
      Benzo_b_fluoranthene:matix = "SED" ;
      Benzo_b_fluoranthene:units = "nanograms/gram" ;
      Benzo_b_fluoranthene:_FillValue = -1. ;
      Benzo_b_fluoranthene:valid_min = 0. ;
      Benzo_b_fluoranthene:valid_max = 1.79769313486232e+308 ;
      Benzo_b_fluoranthene:instrument = "PAH_2002_Sample_dry_weight" ;
      Benzo_b_fluoranthene:grid_mapping = "crs" ;
      Benzo_b_fluoranthene:reference = "0074376/data/0-data/Bioeffects_Assessments/Kachemak_Bay/Data_Files/KB1_ORG.txt" ;
   double Benzo_e_pyrene(Sample_Site) ;
      Benzo_e_pyrene:long_name = "Benzo[e]pyrene" ;
      Benzo_e_pyrene:coordinates = "latitude longitude time z" ;
      Benzo_e_pyrene:matix = "SED" ;
      Benzo_e_pyrene:units = "nanograms/gram" ;
      Benzo_e_pyrene:_FillValue = -1. ;
      Benzo_e_pyrene:valid_min = 0. ;
      Benzo_e_pyrene:valid_max = 1.79769313486232e+308 ;
      Benzo_e_pyrene:instrument = "PAH_2002_Sample_dry_weight" ;
      Benzo_e_pyrene:grid_mapping = "crs" ;
      Benzo_e_pyrene:reference = "0074376/data/0-data/Bioeffects_Assessments/Kachemak_Bay/Data_Files/KB1_ORG.txt" ;
   double Benzo_g_h_i_perylene(Sample_Site) ;
      Benzo_g_h_i_perylene:long_name = "Benzo[g,h,i]perylene" ;
      Benzo_g_h_i_perylene:coordinates = "latitude longitude time z" ;
      Benzo_g_h_i_perylene:matix = "SED" ;
      Benzo_g_h_i_perylene:units = "nanograms/gram" ;
      Benzo_g_h_i_perylene:_FillValue = -1. ;
      Benzo_g_h_i_perylene:valid_min = 0. ;
      Benzo_g_h_i_perylene:valid_max = 1.79769313486232e+308 ;
      Benzo_g_h_i_perylene:instrument = "PAH_2002_Sample_dry_weight" ;
      Benzo_g_h_i_perylene:grid_mapping = "crs" ;
      Benzo_g_h_i_perylene:reference = "0074376/data/0-data/Bioeffects_Assessments/Kachemak_Bay/Data_Files/KB1_ORG.txt" ;
   double Benzo_k_fluoranthene(Sample_Site) ;
      Benzo_k_fluoranthene:long_name = "Benzo[k]fluoranthene" ;
      Benzo_k_fluoranthene:coordinates = "latitude longitude time z" ;
      Benzo_k_fluoranthene:matix = "SED" ;
      Benzo_k_fluoranthene:units = "nanograms/gram" ;
      Benzo_k_fluoranthene:_FillValue = -1. ;
      Benzo_k_fluoranthene:valid_min = 0. ;
      Benzo_k_fluoranthene:valid_max = 1.79769313486232e+308 ;
      Benzo_k_fluoranthene:instrument = "PAH_2002_Sample_dry_weight" ;
      Benzo_k_fluoranthene:grid_mapping = "crs" ;
      Benzo_k_fluoranthene:reference = "0074376/data/0-data/Bioeffects_Assessments/Kachemak_Bay/Data_Files/KB1_ORG.txt" ;
   double Benzothiophene(Sample_Site) ;
      Benzothiophene:long_name = "Benzothiophene" ;
      Benzothiophene:coordinates = "latitude longitude time z" ;
      Benzothiophene:matix = "SED" ;
      Benzothiophene:units = "nanograms/gram" ;
      Benzothiophene:_FillValue = -1. ;
      Benzothiophene:valid_min = 0. ;
      Benzothiophene:valid_max = 1.79769313486232e+308 ;
      Benzothiophene:instrument = "PAH_2002_Sample_dry_weight" ;
      Benzothiophene:grid_mapping = "crs" ;
      Benzothiophene:reference = "0074376/data/0-data/Bioeffects_Assessments/Kachemak_Bay/Data_Files/KB1_ORG.txt" ;
   double Biphenyl(Sample_Site) ;
      Biphenyl:long_name = "Biphenyl" ;
      Biphenyl:coordinates = "latitude longitude time z" ;
      Biphenyl:matix = "SED" ;
      Biphenyl:units = "nanograms/gram" ;
      Biphenyl:_FillValue = -1. ;
      Biphenyl:valid_min = 0. ;
      Biphenyl:valid_max = 1.79769313486232e+308 ;
      Biphenyl:instrument = "PAH_2002_Sample_dry_weight" ;
      Biphenyl:grid_mapping = "crs" ;
      Biphenyl:reference = "0074376/data/0-data/Bioeffects_Assessments/Kachemak_Bay/Data_Files/KB1_ORG.txt" ;
   double C1_Benzothiophene(Sample_Site) ;
      C1_Benzothiophene:long_name = "C1-Benzothiophene" ;
      C1_Benzothiophene:coordinates = "latitude longitude time z" ;
      C1_Benzothiophene:matix = "SED" ;
      C1_Benzothiophene:units = "nanograms/gram" ;
      C1_Benzothiophene:_FillValue = -1. ;
      C1_Benzothiophene:valid_min = 0. ;
      C1_Benzothiophene:valid_max = 1.79769313486232e+308 ;
      C1_Benzothiophene:instrument = "PAH_2002_Sample_dry_weight" ;
      C1_Benzothiophene:grid_mapping = "crs" ;
      C1_Benzothiophene:reference = "0074376/data/0-data/Bioeffects_Assessments/Kachemak_Bay/Data_Files/KB1_ORG.txt" ;
   double C1_Chrysenes(Sample_Site) ;
      C1_Chrysenes:long_name = "C1-Chrysenes" ;
      C1_Chrysenes:coordinates = "latitude longitude time z" ;
      C1_Chrysenes:matix = "SED" ;
      C1_Chrysenes:units = "nanograms/gram" ;
      C1_Chrysenes:_FillValue = -1. ;
      C1_Chrysenes:valid_min = 0. ;
      C1_Chrysenes:valid_max = 1.79769313486232e+308 ;
      C1_Chrysenes:instrument = "PAH_2002_Sample_dry_weight" ;
      C1_Chrysenes:grid_mapping = "crs" ;
      C1_Chrysenes:reference = "0074376/data/0-data/Bioeffects_Assessments/Kachemak_Bay/Data_Files/KB1_ORG.txt" ;
   double C1_Decalin(Sample_Site) ;
      C1_Decalin:long_name = "C1-Decalin" ;
      C1_Decalin:coordinates = "latitude longitude time z" ;
      C1_Decalin:matix = "SED" ;
      C1_Decalin:units = "nanograms/gram" ;
      C1_Decalin:_FillValue = -1. ;
      C1_Decalin:valid_min = 0. ;
      C1_Decalin:valid_max = 1.79769313486232e+308 ;
      C1_Decalin:instrument = "PAH_2002_Sample_dry_weight" ;
      C1_Decalin:grid_mapping = "crs" ;
      C1_Decalin:reference = "0074376/data/0-data/Bioeffects_Assessments/Kachemak_Bay/Data_Files/KB1_ORG.txt" ;
   double C1_Dibenzo_a_h_anthracene(Sample_Site) ;
      C1_Dibenzo_a_h_anthracene:long_name = "C1-Dibenzo[a,h]anthracene" ;
      C1_Dibenzo_a_h_anthracene:coordinates = "latitude longitude time z" ;
      C1_Dibenzo_a_h_anthracene:matix = "SED" ;
      C1_Dibenzo_a_h_anthracene:units = "nanograms/gram" ;
      C1_Dibenzo_a_h_anthracene:_FillValue = -1. ;
      C1_Dibenzo_a_h_anthracene:valid_min = 0. ;
      C1_Dibenzo_a_h_anthracene:valid_max = 1.79769313486232e+308 ;
      C1_Dibenzo_a_h_anthracene:instrument = "PAH_2002_Sample_dry_weight" ;
      C1_Dibenzo_a_h_anthracene:grid_mapping = "crs" ;
      C1_Dibenzo_a_h_anthracene:reference = "0074376/data/0-data/Bioeffects_Assessments/Kachemak_Bay/Data_Files/KB1_ORG.txt" ;
   double C1_Dibenzothiophenes(Sample_Site) ;
      C1_Dibenzothiophenes:long_name = "C1-Dibenzothiophenes" ;
      C1_Dibenzothiophenes:coordinates = "latitude longitude time z" ;
      C1_Dibenzothiophenes:matix = "SED" ;
      C1_Dibenzothiophenes:units = "nanograms/gram" ;
      C1_Dibenzothiophenes:_FillValue = -1. ;
      C1_Dibenzothiophenes:valid_min = 0. ;
      C1_Dibenzothiophenes:valid_max = 1.79769313486232e+308 ;
      C1_Dibenzothiophenes:instrument = "PAH_2002_Sample_dry_weight" ;
      C1_Dibenzothiophenes:grid_mapping = "crs" ;
      C1_Dibenzothiophenes:reference = "0074376/data/0-data/Bioeffects_Assessments/Kachemak_Bay/Data_Files/KB1_ORG.txt" ;
   double C1_Fluoranthenes_Pyrenes(Sample_Site) ;
      C1_Fluoranthenes_Pyrenes:long_name = "C1-Fluoranthenes_Pyrenes" ;
      C1_Fluoranthenes_Pyrenes:coordinates = "latitude longitude time z" ;
      C1_Fluoranthenes_Pyrenes:matix = "SED" ;
      C1_Fluoranthenes_Pyrenes:units = "nanograms/gram" ;
      C1_Fluoranthenes_Pyrenes:_FillValue = -1. ;
      C1_Fluoranthenes_Pyrenes:valid_min = 0. ;
      C1_Fluoranthenes_Pyrenes:valid_max = 1.79769313486232e+308 ;
      C1_Fluoranthenes_Pyrenes:instrument = "PAH_2002_Sample_dry_weight" ;
      C1_Fluoranthenes_Pyrenes:grid_mapping = "crs" ;
      C1_Fluoranthenes_Pyrenes:reference = "0074376/data/0-data/Bioeffects_Assessments/Kachemak_Bay/Data_Files/KB1_ORG.txt" ;
   double C1_Fluorenes(Sample_Site) ;
      C1_Fluorenes:long_name = "C1-Fluorenes" ;
      C1_Fluorenes:coordinates = "latitude longitude time z" ;
      C1_Fluorenes:matix = "SED" ;
      C1_Fluorenes:units = "nanograms/gram" ;
      C1_Fluorenes:_FillValue = -1. ;
      C1_Fluorenes:valid_min = 0. ;
      C1_Fluorenes:valid_max = 1.79769313486232e+308 ;
      C1_Fluorenes:instrument = "PAH_2002_Sample_dry_weight" ;
      C1_Fluorenes:grid_mapping = "crs" ;
      C1_Fluorenes:reference = "0074376/data/0-data/Bioeffects_Assessments/Kachemak_Bay/Data_Files/KB1_ORG.txt" ;
   double C1_Naphthalenes(Sample_Site) ;
      C1_Naphthalenes:long_name = "C1-Naphthalenes" ;
      C1_Naphthalenes:coordinates = "latitude longitude time z" ;
      C1_Naphthalenes:matix = "SED" ;
      C1_Naphthalenes:units = "nanograms/gram" ;
      C1_Naphthalenes:_FillValue = -1. ;
      C1_Naphthalenes:valid_min = 0. ;
      C1_Naphthalenes:valid_max = 1.79769313486232e+308 ;
      C1_Naphthalenes:instrument = "PAH_2002_Sample_dry_weight" ;
      C1_Naphthalenes:grid_mapping = "crs" ;
      C1_Naphthalenes:reference = "0074376/data/0-data/Bioeffects_Assessments/Kachemak_Bay/Data_Files/KB1_ORG.txt" ;
   double C1_Naphthobenzothiophene(Sample_Site) ;
      C1_Naphthobenzothiophene:long_name = "C1-Naphthobenzothiophene" ;
      C1_Naphthobenzothiophene:coordinates = "latitude longitude time z" ;
      C1_Naphthobenzothiophene:matix = "SED" ;
      C1_Naphthobenzothiophene:units = "nanograms/gram" ;
      C1_Naphthobenzothiophene:_FillValue = -1. ;
      C1_Naphthobenzothiophene:valid_min = 0. ;
      C1_Naphthobenzothiophene:valid_max = 1.79769313486232e+308 ;
      C1_Naphthobenzothiophene:instrument = "PAH_2002_Sample_dry_weight" ;
      C1_Naphthobenzothiophene:grid_mapping = "crs" ;
      C1_Naphthobenzothiophene:reference = "0074376/data/0-data/Bioeffects_Assessments/Kachemak_Bay/Data_Files/KB1_ORG.txt" ;
   double C1_Phenanthrenes_Anthracenes(Sample_Site) ;
      C1_Phenanthrenes_Anthracenes:long_name = "C1-Phenanthrenes_Anthracenes" ;
      C1_Phenanthrenes_Anthracenes:coordinates = "latitude longitude time z" ;
      C1_Phenanthrenes_Anthracenes:matix = "SED" ;
      C1_Phenanthrenes_Anthracenes:units = "nanograms/gram" ;
      C1_Phenanthrenes_Anthracenes:_FillValue = -1. ;
      C1_Phenanthrenes_Anthracenes:valid_min = 0. ;
      C1_Phenanthrenes_Anthracenes:valid_max = 1.79769313486232e+308 ;
      C1_Phenanthrenes_Anthracenes:instrument = "PAH_2002_Sample_dry_weight" ;
      C1_Phenanthrenes_Anthracenes:grid_mapping = "crs" ;
      C1_Phenanthrenes_Anthracenes:reference = "0074376/data/0-data/Bioeffects_Assessments/Kachemak_Bay/Data_Files/KB1_ORG.txt" ;
   double C2_Benzothiophene(Sample_Site) ;
      C2_Benzothiophene:long_name = "C2-Benzothiophene" ;
      C2_Benzothiophene:coordinates = "latitude longitude time z" ;
      C2_Benzothiophene:matix = "SED" ;
      C2_Benzothiophene:units = "nanograms/gram" ;
      C2_Benzothiophene:_FillValue = -1. ;
      C2_Benzothiophene:valid_min = 0. ;
      C2_Benzothiophene:valid_max = 1.79769313486232e+308 ;
      C2_Benzothiophene:instrument = "PAH_2002_Sample_dry_weight" ;
      C2_Benzothiophene:grid_mapping = "crs" ;
      C2_Benzothiophene:reference = "0074376/data/0-data/Bioeffects_Assessments/Kachemak_Bay/Data_Files/KB1_ORG.txt" ;
   double C2_Chrysenes(Sample_Site) ;
      C2_Chrysenes:long_name = "C2-Chrysenes" ;
      C2_Chrysenes:coordinates = "latitude longitude time z" ;
      C2_Chrysenes:matix = "SED" ;
      C2_Chrysenes:units = "nanograms/gram" ;
      C2_Chrysenes:_FillValue = -1. ;
      C2_Chrysenes:valid_min = 0. ;
      C2_Chrysenes:valid_max = 1.79769313486232e+308 ;
      C2_Chrysenes:instrument = "PAH_2002_Sample_dry_weight" ;
      C2_Chrysenes:grid_mapping = "crs" ;
      C2_Chrysenes:reference = "0074376/data/0-data/Bioeffects_Assessments/Kachemak_Bay/Data_Files/KB1_ORG.txt" ;
   double C2_Decalin(Sample_Site) ;
      C2_Decalin:long_name = "C2-Decalin" ;
      C2_Decalin:coordinates = "latitude longitude time z" ;
      C2_Decalin:matix = "SED" ;
      C2_Decalin:units = "nanograms/gram" ;
      C2_Decalin:_FillValue = -1. ;
      C2_Decalin:valid_min = 0. ;
      C2_Decalin:valid_max = 1.79769313486232e+308 ;
      C2_Decalin:instrument = "PAH_2002_Sample_dry_weight" ;
      C2_Decalin:grid_mapping = "crs" ;
      C2_Decalin:reference = "0074376/data/0-data/Bioeffects_Assessments/Kachemak_Bay/Data_Files/KB1_ORG.txt" ;
   double C2_Dibenzo_a_h_anthracene(Sample_Site) ;
      C2_Dibenzo_a_h_anthracene:long_name = "C2-Dibenzo[a,h]anthracene" ;
      C2_Dibenzo_a_h_anthracene:coordinates = "latitude longitude time z" ;
      C2_Dibenzo_a_h_anthracene:matix = "SED" ;
      C2_Dibenzo_a_h_anthracene:units = "nanograms/gram" ;
      C2_Dibenzo_a_h_anthracene:_FillValue = -1. ;
      C2_Dibenzo_a_h_anthracene:valid_min = 0. ;
      C2_Dibenzo_a_h_anthracene:valid_max = 1.79769313486232e+308 ;
      C2_Dibenzo_a_h_anthracene:instrument = "PAH_2002_Sample_dry_weight" ;
      C2_Dibenzo_a_h_anthracene:grid_mapping = "crs" ;
      C2_Dibenzo_a_h_anthracene:reference = "0074376/data/0-data/Bioeffects_Assessments/Kachemak_Bay/Data_Files/KB1_ORG.txt" ;
   double C2_Dibenzothiophenes(Sample_Site) ;
      C2_Dibenzothiophenes:long_name = "C2-Dibenzothiophenes" ;
      C2_Dibenzothiophenes:coordinates = "latitude longitude time z" ;
      C2_Dibenzothiophenes:matix = "SED" ;
      C2_Dibenzothiophenes:units = "nanograms/gram" ;
      C2_Dibenzothiophenes:_FillValue = -1. ;
      C2_Dibenzothiophenes:valid_min = 0. ;
      C2_Dibenzothiophenes:valid_max = 1.79769313486232e+308 ;
      C2_Dibenzothiophenes:instrument = "PAH_2002_Sample_dry_weight" ;
      C2_Dibenzothiophenes:grid_mapping = "crs" ;
      C2_Dibenzothiophenes:reference = "0074376/data/0-data/Bioeffects_Assessments/Kachemak_Bay/Data_Files/KB1_ORG.txt" ;
   double C2_Fluoranthenes_Pyrenes(Sample_Site) ;
      C2_Fluoranthenes_Pyrenes:long_name = "C2-Fluoranthenes_Pyrenes" ;
      C2_Fluoranthenes_Pyrenes:coordinates = "latitude longitude time z" ;
      C2_Fluoranthenes_Pyrenes:matix = "SED" ;
      C2_Fluoranthenes_Pyrenes:units = "nanograms/gram" ;
      C2_Fluoranthenes_Pyrenes:_FillValue = -1. ;
      C2_Fluoranthenes_Pyrenes:valid_min = 0. ;
      C2_Fluoranthenes_Pyrenes:valid_max = 1.79769313486232e+308 ;
      C2_Fluoranthenes_Pyrenes:instrument = "PAH_2002_Sample_dry_weight" ;
      C2_Fluoranthenes_Pyrenes:grid_mapping = "crs" ;
      C2_Fluoranthenes_Pyrenes:reference = "0074376/data/0-data/Bioeffects_Assessments/Kachemak_Bay/Data_Files/KB1_ORG.txt" ;
   double C2_Fluorenes(Sample_Site) ;
      C2_Fluorenes:long_name = "C2-Fluorenes" ;
      C2_Fluorenes:coordinates = "latitude longitude time z" ;
      C2_Fluorenes:matix = "SED" ;
      C2_Fluorenes:units = "nanograms/gram" ;
      C2_Fluorenes:_FillValue = -1. ;
      C2_Fluorenes:valid_min = 0. ;
      C2_Fluorenes:valid_max = 1.79769313486232e+308 ;
      C2_Fluorenes:instrument = "PAH_2002_Sample_dry_weight" ;
      C2_Fluorenes:grid_mapping = "crs" ;
      C2_Fluorenes:reference = "0074376/data/0-data/Bioeffects_Assessments/Kachemak_Bay/Data_Files/KB1_ORG.txt" ;
   double C2_Naphthalenes(Sample_Site) ;
      C2_Naphthalenes:long_name = "C2-Naphthalenes" ;
      C2_Naphthalenes:coordinates = "latitude longitude time z" ;
      C2_Naphthalenes:matix = "SED" ;
      C2_Naphthalenes:units = "nanograms/gram" ;
      C2_Naphthalenes:_FillValue = -1. ;
      C2_Naphthalenes:valid_min = 0. ;
      C2_Naphthalenes:valid_max = 1.79769313486232e+308 ;
      C2_Naphthalenes:instrument = "PAH_2002_Sample_dry_weight" ;
      C2_Naphthalenes:grid_mapping = "crs" ;
      C2_Naphthalenes:reference = "0074376/data/0-data/Bioeffects_Assessments/Kachemak_Bay/Data_Files/KB1_ORG.txt" ;
   double C2_Naphthobenzothiophene(Sample_Site) ;
      C2_Naphthobenzothiophene:long_name = "C2-Naphthobenzothiophene" ;
      C2_Naphthobenzothiophene:coordinates = "latitude longitude time z" ;
      C2_Naphthobenzothiophene:matix = "SED" ;
      C2_Naphthobenzothiophene:units = "nanograms/gram" ;
      C2_Naphthobenzothiophene:_FillValue = -1. ;
      C2_Naphthobenzothiophene:valid_min = 0. ;
      C2_Naphthobenzothiophene:valid_max = 1.79769313486232e+308 ;
      C2_Naphthobenzothiophene:instrument = "PAH_2002_Sample_dry_weight" ;
      C2_Naphthobenzothiophene:grid_mapping = "crs" ;
      C2_Naphthobenzothiophene:reference = "0074376/data/0-data/Bioeffects_Assessments/Kachemak_Bay/Data_Files/KB1_ORG.txt" ;
   double C2_Phenanthrenes_Anthracenes(Sample_Site) ;
      C2_Phenanthrenes_Anthracenes:long_name = "C2-Phenanthrenes_Anthracenes" ;
      C2_Phenanthrenes_Anthracenes:coordinates = "latitude longitude time z" ;
      C2_Phenanthrenes_Anthracenes:matix = "SED" ;
      C2_Phenanthrenes_Anthracenes:units = "nanograms/gram" ;
      C2_Phenanthrenes_Anthracenes:_FillValue = -1. ;
      C2_Phenanthrenes_Anthracenes:valid_min = 0. ;
      C2_Phenanthrenes_Anthracenes:valid_max = 1.79769313486232e+308 ;
      C2_Phenanthrenes_Anthracenes:instrument = "PAH_2002_Sample_dry_weight" ;
      C2_Phenanthrenes_Anthracenes:grid_mapping = "crs" ;
      C2_Phenanthrenes_Anthracenes:reference = "0074376/data/0-data/Bioeffects_Assessments/Kachemak_Bay/Data_Files/KB1_ORG.txt" ;
   double C3_Benzothiophene(Sample_Site) ;
      C3_Benzothiophene:long_name = "C3-Benzothiophene" ;
      C3_Benzothiophene:coordinates = "latitude longitude time z" ;
      C3_Benzothiophene:matix = "SED" ;
      C3_Benzothiophene:units = "nanograms/gram" ;
      C3_Benzothiophene:_FillValue = -1. ;
      C3_Benzothiophene:valid_min = 0. ;
      C3_Benzothiophene:valid_max = 1.79769313486232e+308 ;
      C3_Benzothiophene:instrument = "PAH_2002_Sample_dry_weight" ;
      C3_Benzothiophene:grid_mapping = "crs" ;
      C3_Benzothiophene:reference = "0074376/data/0-data/Bioeffects_Assessments/Kachemak_Bay/Data_Files/KB1_ORG.txt" ;
   double C3_Chrysenes(Sample_Site) ;
      C3_Chrysenes:long_name = "C3-Chrysenes" ;
      C3_Chrysenes:coordinates = "latitude longitude time z" ;
      C3_Chrysenes:matix = "SED" ;
      C3_Chrysenes:units = "nanograms/gram" ;
      C3_Chrysenes:_FillValue = -1. ;
      C3_Chrysenes:valid_min = 0. ;
      C3_Chrysenes:valid_max = 1.79769313486232e+308 ;
      C3_Chrysenes:instrument = "PAH_2002_Sample_dry_weight" ;
      C3_Chrysenes:grid_mapping = "crs" ;
      C3_Chrysenes:reference = "0074376/data/0-data/Bioeffects_Assessments/Kachemak_Bay/Data_Files/KB1_ORG.txt" ;
   double C3_Decalin(Sample_Site) ;
      C3_Decalin:long_name = "C3-Decalin" ;
      C3_Decalin:coordinates = "latitude longitude time z" ;
      C3_Decalin:matix = "SED" ;
      C3_Decalin:units = "nanograms/gram" ;
      C3_Decalin:_FillValue = -1. ;
      C3_Decalin:valid_min = 0. ;
      C3_Decalin:valid_max = 1.79769313486232e+308 ;
      C3_Decalin:instrument = "PAH_2002_Sample_dry_weight" ;
      C3_Decalin:grid_mapping = "crs" ;
      C3_Decalin:reference = "0074376/data/0-data/Bioeffects_Assessments/Kachemak_Bay/Data_Files/KB1_ORG.txt" ;
   double C3_Dibenzo_a_h_anthracene(Sample_Site) ;
      C3_Dibenzo_a_h_anthracene:long_name = "C3-Dibenzo[a,h]anthracene" ;
      C3_Dibenzo_a_h_anthracene:coordinates = "latitude longitude time z" ;
      C3_Dibenzo_a_h_anthracene:matix = "SED" ;
      C3_Dibenzo_a_h_anthracene:units = "nanograms/gram" ;
      C3_Dibenzo_a_h_anthracene:_FillValue = -1. ;
      C3_Dibenzo_a_h_anthracene:valid_min = 0. ;
      C3_Dibenzo_a_h_anthracene:valid_max = 1.79769313486232e+308 ;
      C3_Dibenzo_a_h_anthracene:instrument = "PAH_2002_Sample_dry_weight" ;
      C3_Dibenzo_a_h_anthracene:grid_mapping = "crs" ;
      C3_Dibenzo_a_h_anthracene:reference = "0074376/data/0-data/Bioeffects_Assessments/Kachemak_Bay/Data_Files/KB1_ORG.txt" ;
   double C3_Dibenzothiophenes(Sample_Site) ;
      C3_Dibenzothiophenes:long_name = "C3-Dibenzothiophenes" ;
      C3_Dibenzothiophenes:coordinates = "latitude longitude time z" ;
      C3_Dibenzothiophenes:matix = "SED" ;
      C3_Dibenzothiophenes:units = "nanograms/gram" ;
      C3_Dibenzothiophenes:_FillValue = -1. ;
      C3_Dibenzothiophenes:valid_min = 0. ;
      C3_Dibenzothiophenes:valid_max = 1.79769313486232e+308 ;
      C3_Dibenzothiophenes:instrument = "PAH_2002_Sample_dry_weight" ;
      C3_Dibenzothiophenes:grid_mapping = "crs" ;
      C3_Dibenzothiophenes:reference = "0074376/data/0-data/Bioeffects_Assessments/Kachemak_Bay/Data_Files/KB1_ORG.txt" ;
   double C3_Fluoranthenes_Pyrenes(Sample_Site) ;
      C3_Fluoranthenes_Pyrenes:long_name = "C3-Fluoranthenes_Pyrenes" ;
      C3_Fluoranthenes_Pyrenes:coordinates = "latitude longitude time z" ;
      C3_Fluoranthenes_Pyrenes:matix = "SED" ;
      C3_Fluoranthenes_Pyrenes:units = "nanograms/gram" ;
      C3_Fluoranthenes_Pyrenes:_FillValue = -1. ;
      C3_Fluoranthenes_Pyrenes:valid_min = 0. ;
      C3_Fluoranthenes_Pyrenes:valid_max = 1.79769313486232e+308 ;
      C3_Fluoranthenes_Pyrenes:instrument = "PAH_2002_Sample_dry_weight" ;
      C3_Fluoranthenes_Pyrenes:grid_mapping = "crs" ;
      C3_Fluoranthenes_Pyrenes:reference = "0074376/data/0-data/Bioeffects_Assessments/Kachemak_Bay/Data_Files/KB1_ORG.txt" ;
   double C3_Fluorenes(Sample_Site) ;
      C3_Fluorenes:long_name = "C3-Fluorenes" ;
      C3_Fluorenes:coordinates = "latitude longitude time z" ;
      C3_Fluorenes:matix = "SED" ;
      C3_Fluorenes:units = "nanograms/gram" ;
      C3_Fluorenes:_FillValue = -1. ;
      C3_Fluorenes:valid_min = 0. ;
      C3_Fluorenes:valid_max = 1.79769313486232e+308 ;
      C3_Fluorenes:instrument = "PAH_2002_Sample_dry_weight" ;
      C3_Fluorenes:grid_mapping = "crs" ;
      C3_Fluorenes:reference = "0074376/data/0-data/Bioeffects_Assessments/Kachemak_Bay/Data_Files/KB1_ORG.txt" ;
   double C3_Naphthalenes(Sample_Site) ;
      C3_Naphthalenes:long_name = "C3-Naphthalenes" ;
      C3_Naphthalenes:coordinates = "latitude longitude time z" ;
      C3_Naphthalenes:matix = "SED" ;
      C3_Naphthalenes:units = "nanograms/gram" ;
      C3_Naphthalenes:_FillValue = -1. ;
      C3_Naphthalenes:valid_min = 0. ;
      C3_Naphthalenes:valid_max = 1.79769313486232e+308 ;
      C3_Naphthalenes:instrument = "PAH_2002_Sample_dry_weight" ;
      C3_Naphthalenes:grid_mapping = "crs" ;
      C3_Naphthalenes:reference = "0074376/data/0-data/Bioeffects_Assessments/Kachemak_Bay/Data_Files/KB1_ORG.txt" ;
   double C3_Naphthobenzothiophene(Sample_Site) ;
      C3_Naphthobenzothiophene:long_name = "C3-Naphthobenzothiophene" ;
      C3_Naphthobenzothiophene:coordinates = "latitude longitude time z" ;
      C3_Naphthobenzothiophene:matix = "SED" ;
      C3_Naphthobenzothiophene:units = "nanograms/gram" ;
      C3_Naphthobenzothiophene:_FillValue = -1. ;
      C3_Naphthobenzothiophene:valid_min = 0. ;
      C3_Naphthobenzothiophene:valid_max = 1.79769313486232e+308 ;
      C3_Naphthobenzothiophene:instrument = "PAH_2002_Sample_dry_weight" ;
      C3_Naphthobenzothiophene:grid_mapping = "crs" ;
      C3_Naphthobenzothiophene:reference = "0074376/data/0-data/Bioeffects_Assessments/Kachemak_Bay/Data_Files/KB1_ORG.txt" ;
   double C3_Phenanthrenes_Anthracenes(Sample_Site) ;
      C3_Phenanthrenes_Anthracenes:long_name = "C3-Phenanthrenes_Anthracenes" ;
      C3_Phenanthrenes_Anthracenes:coordinates = "latitude longitude time z" ;
      C3_Phenanthrenes_Anthracenes:matix = "SED" ;
      C3_Phenanthrenes_Anthracenes:units = "nanograms/gram" ;
      C3_Phenanthrenes_Anthracenes:_FillValue = -1. ;
      C3_Phenanthrenes_Anthracenes:valid_min = 0. ;
      C3_Phenanthrenes_Anthracenes:valid_max = 1.79769313486232e+308 ;
      C3_Phenanthrenes_Anthracenes:instrument = "PAH_2002_Sample_dry_weight" ;
      C3_Phenanthrenes_Anthracenes:grid_mapping = "crs" ;
      C3_Phenanthrenes_Anthracenes:reference = "0074376/data/0-data/Bioeffects_Assessments/Kachemak_Bay/Data_Files/KB1_ORG.txt" ;
   double C4_Chrysenes(Sample_Site) ;
      C4_Chrysenes:long_name = "C4-Chrysenes" ;
      C4_Chrysenes:coordinates = "latitude longitude time z" ;
      C4_Chrysenes:matix = "SED" ;
      C4_Chrysenes:units = "nanograms/gram" ;
      C4_Chrysenes:_FillValue = -1. ;
      C4_Chrysenes:valid_min = 0. ;
      C4_Chrysenes:valid_max = 1.79769313486232e+308 ;
      C4_Chrysenes:instrument = "PAH_2002_Sample_dry_weight" ;
      C4_Chrysenes:grid_mapping = "crs" ;
      C4_Chrysenes:reference = "0074376/data/0-data/Bioeffects_Assessments/Kachemak_Bay/Data_Files/KB1_ORG.txt" ;
   double C4_Decalin(Sample_Site) ;
      C4_Decalin:long_name = "C4-Decalin" ;
      C4_Decalin:coordinates = "latitude longitude time z" ;
      C4_Decalin:matix = "SED" ;
      C4_Decalin:units = "nanograms/gram" ;
      C4_Decalin:_FillValue = -1. ;
      C4_Decalin:valid_min = 0. ;
      C4_Decalin:valid_max = 1.79769313486232e+308 ;
      C4_Decalin:instrument = "PAH_2002_Sample_dry_weight" ;
      C4_Decalin:grid_mapping = "crs" ;
      C4_Decalin:reference = "0074376/data/0-data/Bioeffects_Assessments/Kachemak_Bay/Data_Files/KB1_ORG.txt" ;
   double C4_Naphthalenes(Sample_Site) ;
      C4_Naphthalenes:long_name = "C4-Naphthalenes" ;
      C4_Naphthalenes:coordinates = "latitude longitude time z" ;
      C4_Naphthalenes:matix = "SED" ;
      C4_Naphthalenes:units = "nanograms/gram" ;
      C4_Naphthalenes:_FillValue = -1. ;
      C4_Naphthalenes:valid_min = 0. ;
      C4_Naphthalenes:valid_max = 1.79769313486232e+308 ;
      C4_Naphthalenes:instrument = "PAH_2002_Sample_dry_weight" ;
      C4_Naphthalenes:grid_mapping = "crs" ;
      C4_Naphthalenes:reference = "0074376/data/0-data/Bioeffects_Assessments/Kachemak_Bay/Data_Files/KB1_ORG.txt" ;
   double C4_Phenanthrenes_Anthracenes(Sample_Site) ;
      C4_Phenanthrenes_Anthracenes:long_name = "C4-Phenanthrenes_Anthracenes" ;
      C4_Phenanthrenes_Anthracenes:coordinates = "latitude longitude time z" ;
      C4_Phenanthrenes_Anthracenes:matix = "SED" ;
      C4_Phenanthrenes_Anthracenes:units = "nanograms/gram" ;
      C4_Phenanthrenes_Anthracenes:_FillValue = -1. ;
      C4_Phenanthrenes_Anthracenes:valid_min = 0. ;
      C4_Phenanthrenes_Anthracenes:valid_max = 1.79769313486232e+308 ;
      C4_Phenanthrenes_Anthracenes:instrument = "PAH_2002_Sample_dry_weight" ;
      C4_Phenanthrenes_Anthracenes:grid_mapping = "crs" ;
      C4_Phenanthrenes_Anthracenes:reference = "0074376/data/0-data/Bioeffects_Assessments/Kachemak_Bay/Data_Files/KB1_ORG.txt" ;
   double Chrysene(Sample_Site) ;
      Chrysene:long_name = "Chrysene" ;
      Chrysene:coordinates = "latitude longitude time z" ;
      Chrysene:matix = "SED" ;
      Chrysene:units = "nanograms/gram" ;
      Chrysene:_FillValue = -1. ;
      Chrysene:valid_min = 0. ;
      Chrysene:valid_max = 1.79769313486232e+308 ;
      Chrysene:instrument = "PAH_2002_Sample_dry_weight" ;
      Chrysene:grid_mapping = "crs" ;
      Chrysene:reference = "0074376/data/0-data/Bioeffects_Assessments/Kachemak_Bay/Data_Files/KB1_ORG.txt" ;
   double Decalin(Sample_Site) ;
      Decalin:long_name = "Decalin" ;
      Decalin:coordinates = "latitude longitude time z" ;
      Decalin:matix = "SED" ;
      Decalin:units = "nanograms/gram" ;
      Decalin:_FillValue = -1. ;
      Decalin:valid_min = 0. ;
      Decalin:valid_max = 1.79769313486232e+308 ;
      Decalin:instrument = "PAH_2002_Sample_dry_weight" ;
      Decalin:grid_mapping = "crs" ;
      Decalin:reference = "0074376/data/0-data/Bioeffects_Assessments/Kachemak_Bay/Data_Files/KB1_ORG.txt" ;
   double Dibenzo_a_h_anthracene(Sample_Site) ;
      Dibenzo_a_h_anthracene:long_name = "Dibenzo[a,h]anthracene" ;
      Dibenzo_a_h_anthracene:coordinates = "latitude longitude time z" ;
      Dibenzo_a_h_anthracene:matix = "SED" ;
      Dibenzo_a_h_anthracene:units = "nanograms/gram" ;
      Dibenzo_a_h_anthracene:_FillValue = -1. ;
      Dibenzo_a_h_anthracene:valid_min = 0. ;
      Dibenzo_a_h_anthracene:valid_max = 1.79769313486232e+308 ;
      Dibenzo_a_h_anthracene:instrument = "PAH_2002_Sample_dry_weight" ;
      Dibenzo_a_h_anthracene:grid_mapping = "crs" ;
      Dibenzo_a_h_anthracene:reference = "0074376/data/0-data/Bioeffects_Assessments/Kachemak_Bay/Data_Files/KB1_ORG.txt" ;
   double Dibenzofuran(Sample_Site) ;
      Dibenzofuran:long_name = "Dibenzofuran" ;
      Dibenzofuran:coordinates = "latitude longitude time z" ;
      Dibenzofuran:matix = "SED" ;
      Dibenzofuran:units = "nanograms/gram" ;
      Dibenzofuran:_FillValue = -1. ;
      Dibenzofuran:valid_min = 0. ;
      Dibenzofuran:valid_max = 1.79769313486232e+308 ;
      Dibenzofuran:instrument = "PAH_2002_Sample_dry_weight" ;
      Dibenzofuran:grid_mapping = "crs" ;
      Dibenzofuran:reference = "0074376/data/0-data/Bioeffects_Assessments/Kachemak_Bay/Data_Files/KB1_ORG.txt" ;
   double Dibenzothiophene(Sample_Site) ;
      Dibenzothiophene:long_name = "Dibenzothiophene" ;
      Dibenzothiophene:coordinates = "latitude longitude time z" ;
      Dibenzothiophene:matix = "SED" ;
      Dibenzothiophene:units = "nanograms/gram" ;
      Dibenzothiophene:_FillValue = -1. ;
      Dibenzothiophene:valid_min = 0. ;
      Dibenzothiophene:valid_max = 1.79769313486232e+308 ;
      Dibenzothiophene:instrument = "PAH_2002_Sample_dry_weight" ;
      Dibenzothiophene:grid_mapping = "crs" ;
      Dibenzothiophene:reference = "0074376/data/0-data/Bioeffects_Assessments/Kachemak_Bay/Data_Files/KB1_ORG.txt" ;
   double Fluoranthene(Sample_Site) ;
      Fluoranthene:long_name = "Fluoranthene" ;
      Fluoranthene:coordinates = "latitude longitude time z" ;
      Fluoranthene:matix = "SED" ;
      Fluoranthene:units = "nanograms/gram" ;
      Fluoranthene:_FillValue = -1. ;
      Fluoranthene:valid_min = 0. ;
      Fluoranthene:valid_max = 1.79769313486232e+308 ;
      Fluoranthene:instrument = "PAH_2002_Sample_dry_weight" ;
      Fluoranthene:grid_mapping = "crs" ;
      Fluoranthene:reference = "0074376/data/0-data/Bioeffects_Assessments/Kachemak_Bay/Data_Files/KB1_ORG.txt" ;
   double Fluorene(Sample_Site) ;
      Fluorene:long_name = "Fluorene" ;
      Fluorene:coordinates = "latitude longitude time z" ;
      Fluorene:matix = "SED" ;
      Fluorene:units = "nanograms/gram" ;
      Fluorene:_FillValue = -1. ;
      Fluorene:valid_min = 0. ;
      Fluorene:valid_max = 1.79769313486232e+308 ;
      Fluorene:instrument = "PAH_2002_Sample_dry_weight" ;
      Fluorene:grid_mapping = "crs" ;
      Fluorene:reference = "0074376/data/0-data/Bioeffects_Assessments/Kachemak_Bay/Data_Files/KB1_ORG.txt" ;
   double Indeno_1_2_3_c_d_pyrene(Sample_Site) ;
      Indeno_1_2_3_c_d_pyrene:long_name = "Indeno[1,2,3-c,d]pyrene" ;
      Indeno_1_2_3_c_d_pyrene:coordinates = "latitude longitude time z" ;
      Indeno_1_2_3_c_d_pyrene:matix = "SED" ;
      Indeno_1_2_3_c_d_pyrene:units = "nanograms/gram" ;
      Indeno_1_2_3_c_d_pyrene:_FillValue = -1. ;
      Indeno_1_2_3_c_d_pyrene:valid_min = 0. ;
      Indeno_1_2_3_c_d_pyrene:valid_max = 1.79769313486232e+308 ;
      Indeno_1_2_3_c_d_pyrene:instrument = "PAH_2002_Sample_dry_weight" ;
      Indeno_1_2_3_c_d_pyrene:grid_mapping = "crs" ;
      Indeno_1_2_3_c_d_pyrene:reference = "0074376/data/0-data/Bioeffects_Assessments/Kachemak_Bay/Data_Files/KB1_ORG.txt" ;
   double Naphthalene(Sample_Site) ;
      Naphthalene:long_name = "Naphthalene" ;
      Naphthalene:coordinates = "latitude longitude time z" ;
      Naphthalene:matix = "SED" ;
      Naphthalene:units = "nanograms/gram" ;
      Naphthalene:_FillValue = -1. ;
      Naphthalene:valid_min = 0. ;
      Naphthalene:valid_max = 1.79769313486232e+308 ;
      Naphthalene:instrument = "PAH_2002_Sample_dry_weight" ;
      Naphthalene:grid_mapping = "crs" ;
      Naphthalene:reference = "0074376/data/0-data/Bioeffects_Assessments/Kachemak_Bay/Data_Files/KB1_ORG.txt" ;
   double Naphthobenzothiophene(Sample_Site) ;
      Naphthobenzothiophene:long_name = "Naphthobenzothiophene" ;
      Naphthobenzothiophene:coordinates = "latitude longitude time z" ;
      Naphthobenzothiophene:matix = "SED" ;
      Naphthobenzothiophene:units = "nanograms/gram" ;
      Naphthobenzothiophene:_FillValue = -1. ;
      Naphthobenzothiophene:valid_min = 0. ;
      Naphthobenzothiophene:valid_max = 1.79769313486232e+308 ;
      Naphthobenzothiophene:instrument = "PAH_2002_Sample_dry_weight" ;
      Naphthobenzothiophene:grid_mapping = "crs" ;
      Naphthobenzothiophene:reference = "0074376/data/0-data/Bioeffects_Assessments/Kachemak_Bay/Data_Files/KB1_ORG.txt" ;
   double Perylene(Sample_Site) ;
      Perylene:long_name = "Perylene" ;
      Perylene:coordinates = "latitude longitude time z" ;
      Perylene:matix = "SED" ;
      Perylene:units = "nanograms/gram" ;
      Perylene:_FillValue = -1. ;
      Perylene:valid_min = 0. ;
      Perylene:valid_max = 1.79769313486232e+308 ;
      Perylene:instrument = "PAH_2002_Sample_dry_weight" ;
      Perylene:grid_mapping = "crs" ;
      Perylene:reference = "0074376/data/0-data/Bioeffects_Assessments/Kachemak_Bay/Data_Files/KB1_ORG.txt" ;
   double Phenanthrene(Sample_Site) ;
      Phenanthrene:long_name = "Phenanthrene" ;
      Phenanthrene:coordinates = "latitude longitude time z" ;
      Phenanthrene:matix = "SED" ;
      Phenanthrene:units = "nanograms/gram" ;
      Phenanthrene:_FillValue = -1. ;
      Phenanthrene:valid_min = 0. ;
      Phenanthrene:valid_max = 1.79769313486232e+308 ;
      Phenanthrene:instrument = "PAH_2002_Sample_dry_weight" ;
      Phenanthrene:grid_mapping = "crs" ;
      Phenanthrene:reference = "0074376/data/0-data/Bioeffects_Assessments/Kachemak_Bay/Data_Files/KB1_ORG.txt" ;
   double Pyrene(Sample_Site) ;
      Pyrene:long_name = "Pyrene" ;
      Pyrene:coordinates = "latitude longitude time z" ;
      Pyrene:matix = "SED" ;
      Pyrene:units = "nanograms/gram" ;
      Pyrene:_FillValue = -1. ;
      Pyrene:valid_min = 0. ;
      Pyrene:valid_max = 1.79769313486232e+308 ;
      Pyrene:instrument = "PAH_2002_Sample_dry_weight" ;
      Pyrene:grid_mapping = "crs" ;
      Pyrene:reference = "0074376/data/0-data/Bioeffects_Assessments/Kachemak_Bay/Data_Files/KB1_ORG.txt" ;
   double PAH_2002_Sample_dry_weight(Sample_Site) ;
      PAH_2002_Sample_dry_weight:long_name = "Sample dry weight" ;
      PAH_2002_Sample_dry_weight:coordinates = "latitude longitude time z" ;
      PAH_2002_Sample_dry_weight:matix = "SED" ;
      PAH_2002_Sample_dry_weight:units = "gram" ;
      PAH_2002_Sample_dry_weight:_FillValue = -1. ;
      PAH_2002_Sample_dry_weight:valid_min = 0. ;
      PAH_2002_Sample_dry_weight:valid_max = 1.79769313486232e+308 ;
      PAH_2002_Sample_dry_weight:instrument = "PAH_2002" ;
      PAH_2002_Sample_dry_weight:grid_mapping = "crs" ;
      PAH_2002_Sample_dry_weight:reference = "0074376/data/0-data/Bioeffects_Assessments/Kachemak_Bay/Data_Files/KB1_ORG.txt" ;
   double PAH_2002_Sample_percent_dry_weight(Sample_Site) ;
      PAH_2002_Sample_percent_dry_weight:long_name = "Sample percent dry weight" ;
      PAH_2002_Sample_percent_dry_weight:coordinates = "latitude longitude time z" ;
      PAH_2002_Sample_percent_dry_weight:matix = "SED" ;
      PAH_2002_Sample_percent_dry_weight:units = "percent" ;
      PAH_2002_Sample_percent_dry_weight:_FillValue = -1. ;
      PAH_2002_Sample_percent_dry_weight:valid_min = 0. ;
      PAH_2002_Sample_percent_dry_weight:valid_max = 100. ;
      PAH_2002_Sample_percent_dry_weight:instrument = "PAH_2002" ;
      PAH_2002_Sample_percent_dry_weight:grid_mapping = "crs" ;
      PAH_2002_Sample_percent_dry_weight:reference = "0074376/data/0-data/Bioeffects_Assessments/Kachemak_Bay/Data_Files/KB1_ORG.txt" ;
   double PAH_2002_Sample_percent_wet_weight(Sample_Site) ;
      PAH_2002_Sample_percent_wet_weight:long_name = "Sample percent wet weight" ;
      PAH_2002_Sample_percent_wet_weight:coordinates = "latitude longitude time z" ;
      PAH_2002_Sample_percent_wet_weight:matix = "SED" ;
      PAH_2002_Sample_percent_wet_weight:units = "percent" ;
      PAH_2002_Sample_percent_wet_weight:_FillValue = -1. ;
      PAH_2002_Sample_percent_wet_weight:valid_min = 0. ;
      PAH_2002_Sample_percent_wet_weight:valid_max = 100. ;
      PAH_2002_Sample_percent_wet_weight:instrument = "PAH_2002" ;
      PAH_2002_Sample_percent_wet_weight:grid_mapping = "crs" ;
      PAH_2002_Sample_percent_wet_weight:reference = "0074376/data/0-data/Bioeffects_Assessments/Kachemak_Bay/Data_Files/KB1_ORG.txt" ;
   double PAH_2002_Sample_wet_weight(Sample_Site) ;
      PAH_2002_Sample_wet_weight:long_name = "Sample wet weight" ;
      PAH_2002_Sample_wet_weight:coordinates = "latitude longitude time z" ;
      PAH_2002_Sample_wet_weight:matix = "SED" ;
      PAH_2002_Sample_wet_weight:units = "gram" ;
      PAH_2002_Sample_wet_weight:_FillValue = -1. ;
      PAH_2002_Sample_wet_weight:valid_min = 0. ;
      PAH_2002_Sample_wet_weight:valid_max = 1.79769313486232e+308 ;
      PAH_2002_Sample_wet_weight:instrument = "PAH_2002" ;
      PAH_2002_Sample_wet_weight:grid_mapping = "crs" ;
      PAH_2002_Sample_wet_weight:reference = "0074376/data/0-data/Bioeffects_Assessments/Kachemak_Bay/Data_Files/KB1_ORG.txt" ;
   double Total_Inorganic_Carbon(Sample_Site) ;
      Total_Inorganic_Carbon:long_name = "Total Inorganic Carbon" ;
      Total_Inorganic_Carbon:coordinates = "latitude longitude time z" ;
      Total_Inorganic_Carbon:matix = "SED" ;
      Total_Inorganic_Carbon:units = "percent" ;
      Total_Inorganic_Carbon:_FillValue = -1. ;
      Total_Inorganic_Carbon:valid_min = 0. ;
      Total_Inorganic_Carbon:valid_max = 100. ;
      Total_Inorganic_Carbon:instrument = "SEDMT_TC" ;
      Total_Inorganic_Carbon:grid_mapping = "crs" ;
      Total_Inorganic_Carbon:reference = "0074376/data/0-data/Bioeffects_Assessments/Kachemak_Bay/Data_Files/KB1_ORG.txt" ;
   double Total_Organic_Carbon(Sample_Site) ;
      Total_Organic_Carbon:long_name = "Total Organic Carbon" ;
      Total_Organic_Carbon:coordinates = "latitude longitude time z" ;
      Total_Organic_Carbon:matix = "SED" ;
      Total_Organic_Carbon:units = "percent" ;
      Total_Organic_Carbon:_FillValue = -1. ;
      Total_Organic_Carbon:valid_min = 0. ;
      Total_Organic_Carbon:valid_max = 100. ;
      Total_Organic_Carbon:instrument = "SEDMT_TC" ;
      Total_Organic_Carbon:grid_mapping = "crs" ;
      Total_Organic_Carbon:reference = "0074376/data/0-data/Bioeffects_Assessments/Kachemak_Bay/Data_Files/KB1_ORG.txt" ;
   double AFS_Sample_percent_dry_weight(Sample_Site) ;
      AFS_Sample_percent_dry_weight:long_name = "Sample percent dry weight" ;
      AFS_Sample_percent_dry_weight:coordinates = "latitude longitude time z" ;
      AFS_Sample_percent_dry_weight:matix = "SED" ;
      AFS_Sample_percent_dry_weight:units = "percent" ;
      AFS_Sample_percent_dry_weight:_FillValue = -1. ;
      AFS_Sample_percent_dry_weight:valid_min = 0. ;
      AFS_Sample_percent_dry_weight:valid_max = 100. ;
      AFS_Sample_percent_dry_weight:instrument = "AFS" ;
      AFS_Sample_percent_dry_weight:grid_mapping = "crs" ;
      AFS_Sample_percent_dry_weight:reference = "0074376/data/0-data/Bioeffects_Assessments/Kachemak_Bay/Data_Files/KB1_TM.txt" ;
   double AFS_Sample_percent_wet_weight(Sample_Site) ;
      AFS_Sample_percent_wet_weight:long_name = "Sample percent wet weight" ;
      AFS_Sample_percent_wet_weight:coordinates = "latitude longitude time z" ;
      AFS_Sample_percent_wet_weight:matix = "SED" ;
      AFS_Sample_percent_wet_weight:units = "percent" ;
      AFS_Sample_percent_wet_weight:_FillValue = -1. ;
      AFS_Sample_percent_wet_weight:valid_min = 0. ;
      AFS_Sample_percent_wet_weight:valid_max = 100. ;
      AFS_Sample_percent_wet_weight:instrument = "AFS" ;
      AFS_Sample_percent_wet_weight:grid_mapping = "crs" ;
      AFS_Sample_percent_wet_weight:reference = "0074376/data/0-data/Bioeffects_Assessments/Kachemak_Bay/Data_Files/KB1_TM.txt" ;
   double AFS_Sample_wet_weight(Sample_Site) ;
      AFS_Sample_wet_weight:long_name = "Sample wet weight" ;
      AFS_Sample_wet_weight:coordinates = "latitude longitude time z" ;
      AFS_Sample_wet_weight:matix = "SED" ;
      AFS_Sample_wet_weight:units = "gram" ;
      AFS_Sample_wet_weight:_FillValue = -1. ;
      AFS_Sample_wet_weight:valid_min = 0. ;
      AFS_Sample_wet_weight:valid_max = 1.79769313486232e+308 ;
      AFS_Sample_wet_weight:instrument = "AFS" ;
      AFS_Sample_wet_weight:grid_mapping = "crs" ;
      AFS_Sample_wet_weight:reference = "0074376/data/0-data/Bioeffects_Assessments/Kachemak_Bay/Data_Files/KB1_TM.txt" ;
   double Selenium(Sample_Site) ;
      Selenium:long_name = "Selenium" ;
      Selenium:coordinates = "latitude longitude time z" ;
      Selenium:matix = "SED" ;
      Selenium:units = "micrograms/gram" ;
      Selenium:_FillValue = -1. ;
      Selenium:valid_min = 0. ;
      Selenium:valid_max = 1.79769313486232e+308 ;
      Selenium:instrument = "AFS_Sample_dry_weight" ;
      Selenium:grid_mapping = "crs" ;
      Selenium:reference = "0074376/data/0-data/Bioeffects_Assessments/Kachemak_Bay/Data_Files/KB1_TM.txt" ;
   double Mercury(Sample_Site) ;
      Mercury:long_name = "Mercury" ;
      Mercury:coordinates = "latitude longitude time z" ;
      Mercury:matix = "SED" ;
      Mercury:units = "micrograms/gram" ;
      Mercury:_FillValue = -1. ;
      Mercury:valid_min = 0. ;
      Mercury:valid_max = 1.79769313486232e+308 ;
      Mercury:instrument = "CVAAS_Sample_dry_weight" ;
      Mercury:grid_mapping = "crs" ;
      Mercury:reference = "0074376/data/0-data/Bioeffects_Assessments/Kachemak_Bay/Data_Files/KB1_TM.txt" ;
   double CVAAS_Sample_percent_dry_weight(Sample_Site) ;
      CVAAS_Sample_percent_dry_weight:long_name = "Sample percent dry weight" ;
      CVAAS_Sample_percent_dry_weight:coordinates = "latitude longitude time z" ;
      CVAAS_Sample_percent_dry_weight:matix = "SED" ;
      CVAAS_Sample_percent_dry_weight:units = "percent" ;
      CVAAS_Sample_percent_dry_weight:_FillValue = -1. ;
      CVAAS_Sample_percent_dry_weight:valid_min = 0. ;
      CVAAS_Sample_percent_dry_weight:valid_max = 100. ;
      CVAAS_Sample_percent_dry_weight:instrument = "CVAAS" ;
      CVAAS_Sample_percent_dry_weight:grid_mapping = "crs" ;
      CVAAS_Sample_percent_dry_weight:reference = "0074376/data/0-data/Bioeffects_Assessments/Kachemak_Bay/Data_Files/KB1_TM.txt" ;
   double CVAAS_Sample_percent_wet_weight(Sample_Site) ;
      CVAAS_Sample_percent_wet_weight:long_name = "Sample percent wet weight" ;
      CVAAS_Sample_percent_wet_weight:coordinates = "latitude longitude time z" ;
      CVAAS_Sample_percent_wet_weight:matix = "SED" ;
      CVAAS_Sample_percent_wet_weight:units = "percent" ;
      CVAAS_Sample_percent_wet_weight:_FillValue = -1. ;
      CVAAS_Sample_percent_wet_weight:valid_min = 0. ;
      CVAAS_Sample_percent_wet_weight:valid_max = 100. ;
      CVAAS_Sample_percent_wet_weight:instrument = "CVAAS" ;
      CVAAS_Sample_percent_wet_weight:grid_mapping = "crs" ;
      CVAAS_Sample_percent_wet_weight:reference = "0074376/data/0-data/Bioeffects_Assessments/Kachemak_Bay/Data_Files/KB1_TM.txt" ;
   double CVAAS_Sample_wet_weight(Sample_Site) ;
      CVAAS_Sample_wet_weight:long_name = "Sample wet weight" ;
      CVAAS_Sample_wet_weight:coordinates = "latitude longitude time z" ;
      CVAAS_Sample_wet_weight:matix = "SED" ;
      CVAAS_Sample_wet_weight:units = "gram" ;
      CVAAS_Sample_wet_weight:_FillValue = -1. ;
      CVAAS_Sample_wet_weight:valid_min = 0. ;
      CVAAS_Sample_wet_weight:valid_max = 1.79769313486232e+308 ;
      CVAAS_Sample_wet_weight:instrument = "CVAAS" ;
      CVAAS_Sample_wet_weight:grid_mapping = "crs" ;
      CVAAS_Sample_wet_weight:reference = "0074376/data/0-data/Bioeffects_Assessments/Kachemak_Bay/Data_Files/KB1_TM.txt" ;
   double Aluminum(Sample_Site) ;
      Aluminum:long_name = "Aluminum" ;
      Aluminum:coordinates = "latitude longitude time z" ;
      Aluminum:matix = "SED" ;
      Aluminum:units = "micrograms/gram" ;
      Aluminum:_FillValue = -1. ;
      Aluminum:valid_min = 0. ;
      Aluminum:valid_max = 1.79769313486232e+308 ;
      Aluminum:instrument = "ICP_Sample_dry_weight" ;
      Aluminum:grid_mapping = "crs" ;
      Aluminum:reference = "0074376/data/0-data/Bioeffects_Assessments/Kachemak_Bay/Data_Files/KB1_TM.txt" ;
   double Chromium(Sample_Site) ;
      Chromium:long_name = "Chromium" ;
      Chromium:coordinates = "latitude longitude time z" ;
      Chromium:matix = "SED" ;
      Chromium:units = "micrograms/gram" ;
      Chromium:_FillValue = -1. ;
      Chromium:valid_min = 0. ;
      Chromium:valid_max = 1.79769313486232e+308 ;
      Chromium:instrument = "ICP_Sample_dry_weight" ;
      Chromium:grid_mapping = "crs" ;
      Chromium:reference = "0074376/data/0-data/Bioeffects_Assessments/Kachemak_Bay/Data_Files/KB1_TM.txt" ;
   double Copper(Sample_Site) ;
      Copper:long_name = "Copper" ;
      Copper:coordinates = "latitude longitude time z" ;
      Copper:matix = "SED" ;
      Copper:units = "micrograms/gram" ;
      Copper:_FillValue = -1. ;
      Copper:valid_min = 0. ;
      Copper:valid_max = 1.79769313486232e+308 ;
      Copper:instrument = "ICP_Sample_dry_weight" ;
      Copper:grid_mapping = "crs" ;
      Copper:reference = "0074376/data/0-data/Bioeffects_Assessments/Kachemak_Bay/Data_Files/KB1_TM.txt" ;
   double Iron(Sample_Site) ;
      Iron:long_name = "Iron" ;
      Iron:coordinates = "latitude longitude time z" ;
      Iron:matix = "SED" ;
      Iron:units = "micrograms/gram" ;
      Iron:_FillValue = -1. ;
      Iron:valid_min = 0. ;
      Iron:valid_max = 1.79769313486232e+308 ;
      Iron:instrument = "ICP_Sample_dry_weight" ;
      Iron:grid_mapping = "crs" ;
      Iron:reference = "0074376/data/0-data/Bioeffects_Assessments/Kachemak_Bay/Data_Files/KB1_TM.txt" ;
   double Manganese(Sample_Site) ;
      Manganese:long_name = "Manganese" ;
      Manganese:coordinates = "latitude longitude time z" ;
      Manganese:matix = "SED" ;
      Manganese:units = "micrograms/gram" ;
      Manganese:_FillValue = -1. ;
      Manganese:valid_min = 0. ;
      Manganese:valid_max = 1.79769313486232e+308 ;
      Manganese:instrument = "ICP_Sample_dry_weight" ;
      Manganese:grid_mapping = "crs" ;
      Manganese:reference = "0074376/data/0-data/Bioeffects_Assessments/Kachemak_Bay/Data_Files/KB1_TM.txt" ;
   double Nickel(Sample_Site) ;
      Nickel:long_name = "Nickel" ;
      Nickel:coordinates = "latitude longitude time z" ;
      Nickel:matix = "SED" ;
      Nickel:units = "micrograms/gram" ;
      Nickel:_FillValue = -1. ;
      Nickel:valid_min = 0. ;
      Nickel:valid_max = 1.79769313486232e+308 ;
      Nickel:instrument = "ICP_Sample_dry_weight" ;
      Nickel:grid_mapping = "crs" ;
      Nickel:reference = "0074376/data/0-data/Bioeffects_Assessments/Kachemak_Bay/Data_Files/KB1_TM.txt" ;
   double ICP_Sample_percent_dry_weight(Sample_Site) ;
      ICP_Sample_percent_dry_weight:long_name = "Sample percent dry weight" ;
      ICP_Sample_percent_dry_weight:coordinates = "latitude longitude time z" ;
      ICP_Sample_percent_dry_weight:matix = "SED" ;
      ICP_Sample_percent_dry_weight:units = "percent" ;
      ICP_Sample_percent_dry_weight:_FillValue = -1. ;
      ICP_Sample_percent_dry_weight:valid_min = 0. ;
      ICP_Sample_percent_dry_weight:valid_max = 100. ;
      ICP_Sample_percent_dry_weight:instrument = "ICP" ;
      ICP_Sample_percent_dry_weight:grid_mapping = "crs" ;
      ICP_Sample_percent_dry_weight:reference = "0074376/data/0-data/Bioeffects_Assessments/Kachemak_Bay/Data_Files/KB1_TM.txt" ;
   double ICP_Sample_percent_wet_weight(Sample_Site) ;
      ICP_Sample_percent_wet_weight:long_name = "Sample percent wet weight" ;
      ICP_Sample_percent_wet_weight:coordinates = "latitude longitude time z" ;
      ICP_Sample_percent_wet_weight:matix = "SED" ;
      ICP_Sample_percent_wet_weight:units = "percent" ;
      ICP_Sample_percent_wet_weight:_FillValue = -1. ;
      ICP_Sample_percent_wet_weight:valid_min = 0. ;
      ICP_Sample_percent_wet_weight:valid_max = 100. ;
      ICP_Sample_percent_wet_weight:instrument = "ICP" ;
      ICP_Sample_percent_wet_weight:grid_mapping = "crs" ;
      ICP_Sample_percent_wet_weight:reference = "0074376/data/0-data/Bioeffects_Assessments/Kachemak_Bay/Data_Files/KB1_TM.txt" ;
   double ICP_Sample_wet_weight(Sample_Site) ;
      ICP_Sample_wet_weight:long_name = "Sample wet weight" ;
      ICP_Sample_wet_weight:coordinates = "latitude longitude time z" ;
      ICP_Sample_wet_weight:matix = "SED" ;
      ICP_Sample_wet_weight:units = "gram" ;
      ICP_Sample_wet_weight:_FillValue = -1. ;
      ICP_Sample_wet_weight:valid_min = 0. ;
      ICP_Sample_wet_weight:valid_max = 1.79769313486232e+308 ;
      ICP_Sample_wet_weight:instrument = "ICP" ;
      ICP_Sample_wet_weight:grid_mapping = "crs" ;
      ICP_Sample_wet_weight:reference = "0074376/data/0-data/Bioeffects_Assessments/Kachemak_Bay/Data_Files/KB1_TM.txt" ;
   double Silicon(Sample_Site) ;
      Silicon:long_name = "Silicon" ;
      Silicon:coordinates = "latitude longitude time z" ;
      Silicon:matix = "SED" ;
      Silicon:units = "micrograms/gram" ;
      Silicon:_FillValue = -1. ;
      Silicon:valid_min = 0. ;
      Silicon:valid_max = 1.79769313486232e+308 ;
      Silicon:instrument = "ICP_Sample_dry_weight" ;
      Silicon:grid_mapping = "crs" ;
      Silicon:reference = "0074376/data/0-data/Bioeffects_Assessments/Kachemak_Bay/Data_Files/KB1_TM.txt" ;
   double Zinc(Sample_Site) ;
      Zinc:long_name = "Zinc" ;
      Zinc:coordinates = "latitude longitude time z" ;
      Zinc:matix = "SED" ;
      Zinc:units = "micrograms/gram" ;
      Zinc:_FillValue = -1. ;
      Zinc:valid_min = 0. ;
      Zinc:valid_max = 1.79769313486232e+308 ;
      Zinc:instrument = "ICP_Sample_dry_weight" ;
      Zinc:grid_mapping = "crs" ;
      Zinc:reference = "0074376/data/0-data/Bioeffects_Assessments/Kachemak_Bay/Data_Files/KB1_TM.txt" ;
   double Antimony(Sample_Site) ;
      Antimony:long_name = "Antimony" ;
      Antimony:coordinates = "latitude longitude time z" ;
      Antimony:matix = "SED" ;
      Antimony:units = "micrograms/gram" ;
      Antimony:_FillValue = -1. ;
      Antimony:valid_min = 0. ;
      Antimony:valid_max = 1.79769313486232e+308 ;
      Antimony:instrument = "ICP_MS_Sample_dry_weight" ;
      Antimony:grid_mapping = "crs" ;
      Antimony:reference = "0074376/data/0-data/Bioeffects_Assessments/Kachemak_Bay/Data_Files/KB1_TM.txt" ;
   double Arsenic(Sample_Site) ;
      Arsenic:long_name = "Arsenic" ;
      Arsenic:coordinates = "latitude longitude time z" ;
      Arsenic:matix = "SED" ;
      Arsenic:units = "micrograms/gram" ;
      Arsenic:_FillValue = -1. ;
      Arsenic:valid_min = 0. ;
      Arsenic:valid_max = 1.79769313486232e+308 ;
      Arsenic:instrument = "ICP_MS_Sample_dry_weight" ;
      Arsenic:grid_mapping = "crs" ;
      Arsenic:reference = "0074376/data/0-data/Bioeffects_Assessments/Kachemak_Bay/Data_Files/KB1_TM.txt" ;
   double Cadmium(Sample_Site) ;
      Cadmium:long_name = "Cadmium" ;
      Cadmium:coordinates = "latitude longitude time z" ;
      Cadmium:matix = "SED" ;
      Cadmium:units = "micrograms/gram" ;
      Cadmium:_FillValue = -1. ;
      Cadmium:valid_min = 0. ;
      Cadmium:valid_max = 1.79769313486232e+308 ;
      Cadmium:instrument = "ICP_MS_Sample_dry_weight" ;
      Cadmium:grid_mapping = "crs" ;
      Cadmium:reference = "0074376/data/0-data/Bioeffects_Assessments/Kachemak_Bay/Data_Files/KB1_TM.txt" ;
   double Lead(Sample_Site) ;
      Lead:long_name = "Lead" ;
      Lead:coordinates = "latitude longitude time z" ;
      Lead:matix = "SED" ;
      Lead:units = "micrograms/gram" ;
      Lead:_FillValue = -1. ;
      Lead:valid_min = 0. ;
      Lead:valid_max = 1.79769313486232e+308 ;
      Lead:instrument = "ICP_MS_Sample_dry_weight" ;
      Lead:grid_mapping = "crs" ;
      Lead:reference = "0074376/data/0-data/Bioeffects_Assessments/Kachemak_Bay/Data_Files/KB1_TM.txt" ;
   double ICP_MS_Sample_percent_dry_weight(Sample_Site) ;
      ICP_MS_Sample_percent_dry_weight:long_name = "Sample percent dry weight" ;
      ICP_MS_Sample_percent_dry_weight:coordinates = "latitude longitude time z" ;
      ICP_MS_Sample_percent_dry_weight:matix = "SED" ;
      ICP_MS_Sample_percent_dry_weight:units = "percent" ;
      ICP_MS_Sample_percent_dry_weight:_FillValue = -1. ;
      ICP_MS_Sample_percent_dry_weight:valid_min = 0. ;
      ICP_MS_Sample_percent_dry_weight:valid_max = 100. ;
      ICP_MS_Sample_percent_dry_weight:instrument = "ICP_MS" ;
      ICP_MS_Sample_percent_dry_weight:grid_mapping = "crs" ;
      ICP_MS_Sample_percent_dry_weight:reference = "0074376/data/0-data/Bioeffects_Assessments/Kachemak_Bay/Data_Files/KB1_TM.txt" ;
   double ICP_MS_Sample_percent_wet_weight(Sample_Site) ;
      ICP_MS_Sample_percent_wet_weight:long_name = "Sample percent wet weight" ;
      ICP_MS_Sample_percent_wet_weight:coordinates = "latitude longitude time z" ;
      ICP_MS_Sample_percent_wet_weight:matix = "SED" ;
      ICP_MS_Sample_percent_wet_weight:units = "percent" ;
      ICP_MS_Sample_percent_wet_weight:_FillValue = -1. ;
      ICP_MS_Sample_percent_wet_weight:valid_min = 0. ;
      ICP_MS_Sample_percent_wet_weight:valid_max = 100. ;
      ICP_MS_Sample_percent_wet_weight:instrument = "ICP_MS" ;
      ICP_MS_Sample_percent_wet_weight:grid_mapping = "crs" ;
      ICP_MS_Sample_percent_wet_weight:reference = "0074376/data/0-data/Bioeffects_Assessments/Kachemak_Bay/Data_Files/KB1_TM.txt" ;
   double ICP_MS_Sample_wet_weight(Sample_Site) ;
      ICP_MS_Sample_wet_weight:long_name = "Sample wet weight" ;
      ICP_MS_Sample_wet_weight:coordinates = "latitude longitude time z" ;
      ICP_MS_Sample_wet_weight:matix = "SED" ;
      ICP_MS_Sample_wet_weight:units = "gram" ;
      ICP_MS_Sample_wet_weight:_FillValue = -1. ;
      ICP_MS_Sample_wet_weight:valid_min = 0. ;
      ICP_MS_Sample_wet_weight:valid_max = 1.79769313486232e+308 ;
      ICP_MS_Sample_wet_weight:instrument = "ICP_MS" ;
      ICP_MS_Sample_wet_weight:grid_mapping = "crs" ;
      ICP_MS_Sample_wet_weight:reference = "0074376/data/0-data/Bioeffects_Assessments/Kachemak_Bay/Data_Files/KB1_TM.txt" ;
   double Silver(Sample_Site) ;
      Silver:long_name = "Silver" ;
      Silver:coordinates = "latitude longitude time z" ;
      Silver:matix = "SED" ;
      Silver:units = "micrograms/gram" ;
      Silver:_FillValue = -1. ;
      Silver:valid_min = 0. ;
      Silver:valid_max = 1.79769313486232e+308 ;
      Silver:instrument = "ICP_MS_Sample_dry_weight" ;
      Silver:grid_mapping = "crs" ;
      Silver:reference = "0074376/data/0-data/Bioeffects_Assessments/Kachemak_Bay/Data_Files/KB1_TM.txt" ;
   double Tin(Sample_Site) ;
      Tin:long_name = "Tin" ;
      Tin:coordinates = "latitude longitude time z" ;
      Tin:matix = "SED" ;
      Tin:units = "micrograms/gram" ;
      Tin:_FillValue = -1. ;
      Tin:valid_min = 0. ;
      Tin:valid_max = 1.79769313486232e+308 ;
      Tin:instrument = "ICP_MS_Sample_dry_weight" ;
      Tin:grid_mapping = "crs" ;
      Tin:reference = "0074376/data/0-data/Bioeffects_Assessments/Kachemak_Bay/Data_Files/KB1_TM.txt" ;
   double time(Sample_Site) ;
      time:long_name = "time" ;
      time:standard_name = "time" ;
      time:units = "days since 1970-01-01 00:00:00" ;
      time:_FillValue = -1. ;
      time:calendar = "julian" ;
      time:axis = "T" ;
      
   double z(Sample_Site) ;
      z:long_name = "depth below sea level" ;
      z:standard_name = "altitude" ;
      z:units = "meters" ;
      z:positive = "down" ;
      z:_FillValue = -1. ;
      z:axis = "Z" ;
      
   double longitude(Sample_Site) ;
      longitude:long_name = "longitude" ;
      longitude:standard_name = "longitude" ;
      longitude:nodc_name = "longitude" ;
      longitude:units = "degrees_east" ;
      longitude:_FillValue = -999. ;
      longitude:valid_min = -180. ;
      longitude:valid_max = 180. ;
      longitude:axis = "X" ;
      
   double latitude(Sample_Site) ;
      latitude:long_name = "latitude" ;
      latitude:standard_name = "latitude" ;
      latitude:nodc_name = "latitude" ;
      latitude:units = "degrees_north" ;
      latitude:_FillValue = -999. ;
      latitude:valid_min = -90. ;
      latitude:valid_max = 90. ;
      latitude:axis = "Y" ;
      
   char site_code(Sample_Site, NST_Site_code_string_length) ;
      site_code:long_name = "National Status and Trends Program Unique Site Code" ;
      site_code:nodc_name = "Originator_Station_Code" ;
   char site_name(Sample_Site, Site_name_string_length) ;
      site_name:long_name = "Site_Long_Name" ;
   double AFS ;
      AFS:long_name = "" ;
   double AMP_AA ;
      AMP_AA:long_name = "" ;
   double AMP_EE ;
      AMP_EE:long_name = "" ;
   double CVAAS ;
      CVAAS:long_name = "" ;
   double ECDDUAL_M ;
      ECDDUAL_M:long_name = "" ;
   double GS ;
      GS:long_name = "" ;
   double Hexylation ;
      Hexylation:long_name = "" ;
   double ICP ;
      ICP:long_name = "" ;
   double ICP_MS ;
      ICP_MS:long_name = "" ;
   double PAH_2002 ;
      PAH_2002:long_name = "" ;
   double SEDMT_TC ;
      SEDMT_TC:long_name = "" ;
   double crs ;
      crs:grid_mapping_name = "latitude_longitude" ;

// global attributes:
      :title = "Bioeffects Program - Kachemak Bay Database" ;
      :summary = "No summary provided" ;
      :geospatial_lat_min = "59.34" ;
      :geospatial_lat_max = "59.78" ;
      :geospatial_lat_resolution = "~100 meters" ;
      :geospatial_lat_units = "degrees_north" ;
      :geospatial_lon_min = "-151.8" ;
      :geospatial_lon_max = "-151.1" ;
      :geospatial_lon_resolution = "~100 meters" ;
      :geospatial_lon_units = "degrees_east" ;
      :institution = "US DOC; NOAA; NATIONAL OCEAN SERVICE; NATIONAL CENTERS FOR COASTAL OCEAN SCIENCE" ;
      :date_created = "2012-01-30" ;
      :date_modified = "2012-01-30" ;
      :creator_name = "Jonathan N. Blythe, Ph.D." ;
      :creator_url = "www.nodc.noaa.gov" ;
      :contributor_name = "Stuart Ian Hartwell, Oren Perez" ;
      :contributor_role = "Submitter, Producer" ;
      :project = "NATIONAL STATUS and TRENDS" ;
      :keywords = "BENTHIC COMMUNITIES, BIOASSAY, BIOCHEMISTRY, CHEMISTRY - SEDIMENT, METALS, PAH, TRACE METALS" ;
      :keywords_vocabulary = "NODC DATA TYPES THESAURUS" ;
      :references = "NODC Accession 0074376" ;
      :comment = "Laboratory analyses of field collected samples for monitoring marine environmental quality" ;
      :publisher_name = "NOAA/NESDIS/NODC - US National Oceanographic Data Center" ;
      :publisher_email = "NODC.services@noaa.gov" ;
      :publisher_url = "www.nodc.noaa.gov" ;
      :history = "" ;
      :processing_level = "" ;
      :id = "" ;
      :naming_authority = "gov.noaa.nodc" ;
      :license = "none" ;
      :featureType = "station" ;
      :cdm_data_type = "Point" ;
      :nodc_template_version = "NODC_Point_Template_v1.1" ;
      :Conventions = "CF-1.6" ;
      :standard_name_vocabulary = "NetCDF Climate and Forecast (CF) Metadata Convention Standard Name Table v23" ;
      :Metadata_Conventions = "Unidata Dataset Discovery v1.0" ;
      :metadata_link = "0074376/data/0-data/Bioeffects_Assessments/Kachemak_Bay/Metadata/" ;
      :time_coverage_start = "20070810T000000" ;
      :time_coverage_end = "20070814T000000" ;
      :time_coverage_resolution = "day" ;
      :geospatial_vertical_min = 0.9 ;
      :geospatial_vertical_max = 23.8 ;
      :geospatial_vertical_units = "meter" ;
      :geospatial_vertical_positive = "down" ;
}

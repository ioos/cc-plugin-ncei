netcdf NODC_timeseries_orthogonal {
dimensions:
       time = 1;//.................................................... REQUIRED - Number of time steps in the time series
       timeSeries = 2; //............................................... REQUIRED - Number of time series (=1 for single time series or can be removed)
variables:
        int station_id(timeSeries); //....................................... RECOMMENDED - If using the attribute below: cf_role. Data type can be whatever is appropriate for the unique feature type.
                station_id:long_name = "Unique identifier for each feature instance"; //................................ RECOMMENDED
                station_id:cf_role = "timeseries_id"; //..................... RECOMMENDED
        double time(time) ;//........................................ Depending on the precision used for the variable, the data type could be int or double instead of float.
                time:long_name = "Time" ; //..................................... RECOMMENDED - Provide a descriptive, long name for this variable. 
                time:standard_name = "time" ; //............................. REQUIRED    - Do not change
                time:units = "seconds since 1970-01-01T00:00:00Z" ; //... REQUIRED    - Use approved CF convention with approved UDUNITS.
                time:axis = "T" ; //......................................... REQUIRED    - Do not change.
                time:comment = "Time as reported by the controller clock" ; //....................................... RECOMMENDED - Add useful, additional information here.  
        float lat(timeSeries) ;//....................................... Depending on the precision used for the variable, the data type could be int or double instead of float. 
                lat:long_name = "Latitude" ; //...................................... RECOMMENDED - Provide a descriptive, long name for this variable.
                lat:standard_name = "latitude" ; //.......................... REQUIRED    - Do not change.
                lat:units = "degrees_north" ; //............................. REQUIRED    - CF recommends degrees_north, but at least must use UDUNITS.
                lat:axis = "Y" ; //.......................................... REQUIRED    - Do not change.
                lat:valid_min = 41.232f ; //.................................... RECOMMENDED - Replace with correct value.
                lat:valid_max = 41.288f ; //.................................... RECOMMENDED - Replace with correct value.
                lat:comment = "GPS Latitude" ; //........................................ RECOMMENDED - Add useful, additional information here.
       float lon(timeSeries) ; //........................................ Depending on the precision used for the variable, the data type could be int or double instead of float. 
                lon:long_name = "Longitude" ; //...................................... RECOMMENDED
                lon:standard_name = "longitude" ; //......................... REQUIRED    - This is fixed, do not change.
                lon:units = "degrees_east" ; //.............................. REQUIRED    - CF recommends degrees_east, but at least use UDUNITS.
                lon:axis = "X" ; //.......................................... REQUIRED    - Do not change.
                lon:valid_min = -71.772f ; //.................................... RECOMMENDED - Replace this with correct value.
                lon:valid_max = -71.673f ; //.................................... RECOMMENDED - Replace this with correct value.
                lon:comment = "GPS Longitude" ; //........................................ RECOMMENDED - Add useful, additional information here.
        float z(timeSeries) ;//........................................ Depending on the precision used for the variable, the data type could be int or double instead of float. Also the variable "z" could be substituted with a more descriptive name like "depth", "altitude", "pressure", etc.
                z:long_name = "Depth" ; //........................................ RECOMMENDED - Provide a descriptive, long name for this variable. 
                z:standard_name = "depth" ; //.................................... REQUIRED    - Usually "depth" or "altitude" is used.
                z:units = "m" ; //............................................ REQUIRED    - Use UDUNITS.
                z:axis = "Z" ; //............................................ REQUIRED    - Do not change.
                z:positive = "down" ; //......................................... REQUIRED    - Use "up" or "down".
                z:valid_min = 0.0f ; //...................................... RECOMMENDED - Replace with correct value.
                z:valid_max = 0.0f ; //...................................... RECOMMENDED - Replace with correct value.
                z:comment = "Sensors are positioned at water surface" ; //.......................................... RECOMMENDED - Add useful, additional information here.
        float temperature(timeSeries,time) ;//................................ This is an example of how each and every geophysical variable in the file should be represented. Replace the name of the variable("temperature") with a suitable name. Replace "float" by data type which is appropriate for the variable. 
                temperature:long_name = "Temperature" ; //................... RECOMMENDED - Provide a descriptive, long name for this variable. 
                temperature:standard_name = "sea_water_temperature" ; //............... REQUIRED    - If using a CF standard name and a suitable name exists in the CF standard name table.
                temperature:units = "deg_C" ; //....................... REQUIRED    - Use UDUNITS compatible units.
                temperature:_FillValue = -9999.0f ; //................ REQUIRED  if there could be missing values in the data.
                temperature:valid_min = -20.0f ; //................. RECOMMENDED - Replace with correct value.
                temperature:valid_max = 40.0f ; //................. RECOMMENDED - Replace with correct value.
                temperature:coordinates = "time lat lon z" ; //... REQUIRED    - Include the auxiliary coordinate variables and optionally coordinate variables in the list. The order itself does not matter. Also, note that whenever any auxiliary coordinate variable contains a missing value, all other coordinate, auxiliary coordinate and data values corresponding to that element should also contain missing values.
                temperature:grid_mapping = "crs" ; //............. RECOMMENDED - It is highly recommended that the data provider put the data in a well known geographic coordinate system and provide the details of the coordinate system.
                temperature:source = "SBE 37" ; //...................... RECOMMENDED - The method of production of the original data
                temperature:references = "http://www.seabird.com/sbe37si-microcat-ctd" ; //.................. RECOMMENDED - Published or web-based references that describe the data or methods used to produce it.
                temperature: cell_methods = "time: point lon: point lat: point z: point" ; // .............. RECOMMENDED - Use the coordinate variables to define the cell values (ex., "time: point lon: point lat: point z: point").
                temperature:ancillary_variables = "temperature_qc temperature_spike_qc" ; //......... RECOMMENDED - Identify the variable name(s) of the flag(s) and other ancillary variables relevant to this variable.  Use a space-separated list.
                temperature:platform = "platform" ; //... RECOMMENDED - Refers to name of variable containing information on the platform from which this variable was collected.
                temperature:instrument = "instrument_variable";//..RECOMMENDED - Refers to name of variable containing information on the instrument from which this variable was collected.
                temperature:comment = "temperature measured from CTD" ; //..................... RECOMMENDED - Add useful, additional information here.
                temperature:instrument = "ctd_id" ;
        int temperature_qc(timeSeries,time);  //...................... An enumerated flag variable, in which numeric values refer to defined, exclusive conditions.
                temperature_qc:standard_name = "sea_water_temperature status_flag" ; //.............. RECOMMENDED - This attribute should include the standard name of the variable which this flag contributes plus the modifier: "status_flag" (for example, "sea_water_temperature status_flag"). See CF standard name modifiers.
                temperature_qc:long_name = "Temperature Primary QC" ; //................. RECOMMENDED - Provide a descriptive, long name for this variable. 
                temperature_qc:flag_values = 1b, 2b, 3b, 4b, 9b; //.................. REQUIRED    - Provide a comma-separated list of flag values that map to the flag_meanings.
                temperature_qc:flag_meanings = "good not_evaluated suspect bad missing" ; //............. REQUIRED    - Provide a space-separated list of meanings corresponding to each of the flag_values
                temperature_qc:references = "https://ioos.noaa.gov/project/qartod/" ; //................ RECOMMENDED - Published or web-based references that describe the data or methods used to produce it.
                temperature_qc:comment = "Tests performed are global range and spike tests" ; //................... RECOMMENDED - Add useful, additional information here.
        int temperature_spike_qc(timeSeries,time);  //...................... An enumerated flag variable, in which numeric values refer to defined, exclusive conditions.
                temperature_spike_qc:standard_name = "sea_water_temperature status_flag" ; //.............. RECOMMENDED - This attribute should include the standard name of the variable which this flag contributes plus the modifier: "status_flag" (for example, "sea_water_temperature status_flag"). See CF standard name modifiers.
                temperature_spike_qc:long_name = "Temperature Spike QC" ; //................. RECOMMENDED - Provide a descriptive, long name for this variable. 
                temperature_spike_qc:flag_values = 1b, 2b, 3b, 4b, 9b; //.................. REQUIRED    - Provide a comma-separated list of flag values that map to the flag_meanings.
                temperature_spike_qc:flag_meanings = "good not_evaluated suspect bad missing" ; //............. REQUIRED    - Provide a space-separated list of meanings corresponding to each of the flag_values
                temperature_spike_qc:references = "https://ioos.noaa.gov/project/qartod/" ; //................ RECOMMENDED - Published or web-based references that describe the data or methods used to produce it.
                temperature_spike_qc:comment = "Spike test for Temperature" ; //................... RECOMMENDED - Add useful, additional information here.
        int platform; //............................................ RECOMMENDED - a container variable storing information about the platform. If more than one, can expand each attribute into a variable. For example, platform_call_sign and platform_nodc_code. See instrument_parameter_variable for an example.
                platform:long_name = "Coastal Inshore surface platform" ; //........................ RECOMMENDED - Provide a descriptive, long name for this variable. 
                platform:comment = "Equipped with iridium, SBD and GPS" ; //.......................... RECOMMENDED - Add useful, additional information here.
                platform:call_sign = "maverick" ; //........................ RECOMMENDED - This attribute identifies the call sign of the platform. 	 
        int ctd_id; //.................... RECOMMENDED - an instrument variable storing information about a parameter of the instrument used in the measurement, the dimensions don't have to be specified if the same instrument is used for all the measurements.
                ctd_id:long_name = "CTD Identifier" ; //............ RECOMMENDED - Provide a descriptive, long name for this variable. 
                ctd_id:comment = "Each instrument is a CTD SeaBird" ; //.............. RECOMMENDED - Add useful, additional information here.
                ctd_id:serial_numbers = "abc123 321bca" ;
        int crs; //.......................................................... RECOMMENDED - A container variable storing information about the grid_mapping. All the attributes within a grid_mapping variable are described in http://cf-pcmdi.llnl.gov/documents/cf-conventions/1.6/cf-conventions.html#appendix-grid-mappings. For all the measurements based on WSG84, the default coordinate system used for GPS measurements, the values shown here should be used.
                crs:grid_mapping_name = "latitude_longitude"; //............. RECOMMENDED
                crs:epsg_code = "EPSG:4326" ; //............................. RECOMMENDED - European Petroleum Survey Group code for the grid mapping name.
                crs:semi_major_axis = 6378137.0 ; //......................... RECOMMENDED
                crs:inverse_flattening = 298.257223563 ; //.................. RECOMMENDED
// global attributes:
        :Conventions = "CF-1.6" ; //......................................... REQUIRED    - Always try to use latest value. (CF)
        :Metadata_Conventions = "Unidata Dataset Discovery v1.0" ; //........ REQUIRED    - Do not change. (ACDD)
        :featureType = "timeSeries" ; //..................................... REQUIRED - CF attribute for identifying the featureType.
        :cdm_data_type = "Station" ; //...................................... REQUIRED (ACDD)
        :nodc_template_version = "NODC_NetCDF_TimeSeries_Orthogonal_Template_v1.1" ; //....... REQUIRED (NODC)
        :standard_name_vocabulary = "NetCDF Climate and Forecast (CF) Metadata Convention Standard Name Table \"33\"" ; //........ REQUIRED    - If using CF standard name attribute for variables. "X" denotes the table number  (ACDD)
        :title = "Example Multi-station time series" ; //..................................................... RECOMMENDED - Provide a useful title for the data in the file. (ACDD)
        :summary = "Example dataset for the sole purpose of testing the IOOS Compliance Checker" ; //................................................... RECOMMENDED - Provide a useful summary or abstract for the data in the file. (ACDD)
        :source = "raw observations from instruments" ; //.................................................... RECOMMENDED - The input data sources regardless of the method of production method used. (CF)
        :platform = "platform" ; //................................. RECOMMENDED - Refers to a variable containing information about the platform. May also put this in individual variables. Use NODC or ICES platform table. (NODC)
        :uuid = "4e1243bd22c66e76c2ba9eddc1f91394e57f9f83" ; //...................................................... RECOMMENDED - Machine readable unique identifier for each file. A new uuid is created whenever the file is changed. (NODC)
        :sea_name = "Long Island Sound" ; //.................................................. RECOMMENDED - The names of the sea in which the data were collected. Use NODC sea names table. (NODC)
        :id = "Example dataset" ; //........................................................ RECOMMENDED - Should be a human readable unique identifier for data set. (ACDD)
        :naming_authority = "gov.noaa.ioos" ; //.......................................... RECOMMENDED - Backward URL of institution (for example, gov.noaa.nodc). (ACDD)
        :time_coverage_start = "2016-05-22T00:00Z" ; //....................................... RECOMMENDED - Use ISO8601 for date and time. (ACDD)
        :time_coverage_end = "2016-05-23T00:00Z" ; //......................................... RECOMMENDED - Use ISO8601 for date and time.(ACDD)
        :time_coverage_resolution = "hour" ; //.................................. RECOMMENDED - For example, "point" or "minute averages". (ACDD)
        :geospatial_lat_min = 41.232f ; //...................................... RECOMMENDED - Replace with correct value. (ACDD)
        :geospatial_lat_max = 41.288f ; //...................................... RECOMMENDED - Replace with correct value. (ACDD)
        :geospatial_lat_units = "degrees_north" ; //......................... RECOMMENDED - Use UDUNITS compatible units. (ACDD)
        :geospatial_lat_resolution= "point" ; //.................................. RECOMMENDED - For example, "point" or "10 degree grid". (ACDD)
        :geospatial_lon_min = -71.772f ; //...................................... RECOMMENDED - Replace with correct value. (ACDD)
        :geospatial_lon_max = -71.673f ; //...................................... RECOMMENDED - Replace with correct value. (ACDD)
        :geospatial_lon_units = "degrees_east"; //........................... RECOMMENDED - Use UDUNITS compatible units. (ACDD)
        :geospatial_lon_resolution= "point" ; //.................................. RECOMMENDED - For example, "point" or "10 degree grid". (ACDD)
        :geospatial_vertical_min = 0.0f ; //................................. RECOMMENDED - Replace with correct value. (ACDD)
        :geospatial_vertical_max = 0.0f ; //................................. RECOMMENDED - Replace with correct value. (ACDD)
        :geospatial_vertical_units = "m" ; //................................. RECOMMENDED - Use UDUNITS compatible units. (ACDD)
        :geospatial_vertical_resolution = "point" ; //............................ RECOMMENDED - For example, "point" or "1 meter binned". (ACDD)
        :geospatial_vertical_positive = "down" ; //.............................. RECOMMENDED - Use "up" or "down". (ACDD)
        :institution = "NOAA" ; //............................................... RECOMMENDED - Institution of the person or group that collected the data.  An institution attribute can be used for each variable if variables come from more than one institution. (ACDD)
        :creator_name = "Luke Campbell" ; //.............................................. RECOMMENDED - Name of the person who collected the data. (ACDD)
        :creator_url = "https://github.com/lukecampbell/" ; //............................................... RECOMMENDED - URL for person who collected the data. (ACDD)
        :creator_email = "luke.s.campbell-nospam at rpsgroup.com  Remove the -nospam part" ; //............................................. RECOMMENDED - Email address for person who collected the data. (ACDD)
        :project = "IOOS Compliance Checker" ; //................................................... RECOMMENDED - Project the data was collected under. (ACDD)
        :processing_level = "L1" ; //.......................................... RECOMMENDED - Provide a description of the processing or quality control level of the data. (ACDD)
        :references = "https://www.nodc.noaa.gov/data/formats/netcdf/v1.1/timeSeriesOrthogonal.cdl" ; //................................................ RECOMMENDED - Published or web-based references that describe the data or methods used to produce it. (CF)
        :keywords_vocabulary = "Luke" ; //....................................... RECOMMENDED - Identifies the controlled keyword vocabulary used to specify the values within the attribute "keywords". e.g. NASA/GCMD Earth Science Keywords (ACDD)
        :keywords = "Testing" ; //.................................................. RECOMMENDED - A comma separated list of keywords coming from the keywords_vocabulary. (ACDD)
        :acknowledgment = "Testing" ; //............................................ RECOMMENDED - Text to use to properly acknowledge use of the data. (ACDD)
        :comment = "Testing" ; //................................................... RECOMMENDED - Provide useful additional information here. (ACDD and CF)
        :contributor_name = "Testing" ; //.......................................... RECOMMENDED - A comma separated list of contributors to this data set. (ACDD)
        :contributor_role = "Testing" ; //.......................................... RECOMMENDED - A comma separated list of their roles. (ACDD)
        :date_created = "2016-05-23T00:00Z" ; //.............................................. RECOMMENDED - Creation date of the netCDF.  Use ISO8601 for date and time. (ACDD)
        :date_modified = "2016-05-23T00:00Z" ; //............................................. RECOMMENDED - Modification date of the netCDF.  Use ISO8601 for date and time. (ACDD)
        :publisher_name = "Testing" ; //............................................ RECOMMENDED - Publisher of the data. (ACDD)
        :publisher_email = "testing@ioos.us" ; //........................................... RECOMMENDED - Email address of the publisher of the data. (ACDD)
        :publisher_url = "http://ioos.us/" ; //............................................. RECOMMENDED - A URL for the publisher of the data. (ACDD)
        :history = "2016-05-23: Created the file" ; //................................................... RECOMMENDED - Record changes made to the netCDF. (ACDD)
        :license = "Do what you wish, but the data is completely made up and should only be used for testing. And even then it's questionable." ; //................................................... RECOMMENDED - Describe the restrictions to data access and distribution. (ACDD)
        :metadata_link = "http://www.wikipedia.org/" ; //............................................. RECOMMENDED - This attribute provides a link to a complete metadata record for this data set or the collection that contains this data set. (ACDD)    
}

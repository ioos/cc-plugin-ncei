netcdf NCEI_trajectoryProfile_template_v2.0_2016-09-22_181616.896731 {
dimensions:
	obs = 10 ;
	trajectory = 1 ;
	z = 4 ;
variables:
	int trajectory(trajectory) ;
		trajectory:long_name = "Transect 1" ;
		trajectory:cf_role = "trajectory_id" ;
	double time(trajectory, obs) ;
		time:_FillValue = -9999. ;
		time:long_name = "Time" ;
		time:standard_name = "time" ;
		time:units = "seconds since 1970-01-01 00:00:00 UTC" ;
		time:axis = "T" ;
		time:calendar = "julian" ;
		time:comment = "These data are bogus!!!!!" ;
	double lat(trajectory, obs) ;
		lat:_FillValue = -9999. ;
		lat:long_name = "Latitude" ;
		lat:standard_name = "latitude" ;
		lat:units = "degrees_north" ;
		lat:axis = "Y" ;
		lat:valid_min = -90. ;
		lat:valid_max = 90. ;
		lat:comment = "These data are bogus!!!!!" ;
	double lon(trajectory, obs) ;
		lon:_FillValue = -9999. ;
		lon:long_name = "Longitude" ;
		lon:standard_name = "longitude" ;
		lon:units = "degrees_east" ;
		lon:axis = "X" ;
		lon:valid_min = -180. ;
		lon:valid_max = 180. ;
		lon:comment = "These data are bogus!!!!!" ;
	double z(z) ;
		z:long_name = "depth of sensor" ;
		z:standard_name = "depth" ;
		z:units = "m" ;
		z:axis = "Z" ;
		z:valid_min = 0. ;
		z:valid_max = 10971. ;
		z:positive = "down" ;
		z:comment = "These data are bogus!!!!!" ;
	double sal(trajectory, obs, z) ;
		sal:_FillValue = -9999. ;
		sal:long_name = "Salinity" ;
		sal:standard_name = "sea_water_salinity" ;
		sal:units = "0.001" ;
		sal:scale_factor = 1. ;
		sal:add_offset = 0. ;
		sal:valid_min = 0. ;
		sal:valid_max = 100. ;
		sal:data_min = 33.0875659393347 ;
		sal:data_max = 35.9176790819942 ;
		sal:coordinates = "time lat lon z" ;
		sal:coverage_content_type = "physicalMeasurement" ;
		sal:missing_value = -8888. ;
		sal:ncei_name = "SALINITY" ;
		sal:grid_mapping = "crs" ;
		sal:source = "numpy.random.rand function." ;
		sal:references = "http://www.numpy.org/" ;
		sal:cell_methods = "time: point longitude: point latitude: point" ;
		sal:platform = "platform1" ;
		sal:instrument = "instrument1" ;
		sal:comment = "These data are bogus!!!!!" ;
	double temp(trajectory, obs, z) ;
		temp:_FillValue = -9999. ;
		temp:long_name = "Temperature" ;
		temp:standard_name = "sea_water_temperature" ;
		temp:units = "degree_Celsius" ;
		temp:scale_factor = 1. ;
		temp:add_offset = 0. ;
		temp:valid_min = 0. ;
		temp:valid_max = 100. ;
		temp:data_min = 13.1602940932013 ;
		temp:data_max = 15.8440344906993 ;
		temp:coordinates = "time lat lon z" ;
		temp:coverage_content_type = "physicalMeasurement" ;
		temp:missing_value = -8888. ;
		temp:ncei_name = "WATER TEMPERATURE" ;
		temp:grid_mapping = "crs" ;
		temp:source = "numpy.random.rand function." ;
		temp:references = "http://www.numpy.org/" ;
		temp:cell_methods = "time: point longitude: point latitude: point" ;
		temp:platform = "platform1" ;
		temp:instrument = "instrument1" ;
		temp:comment = "These data are bogus!!!!!" ;
	char instrument1 ;
		instrument1:long_name = "Seabird 37 Microcat" ;
		instrument1:ncei_name = "CTD" ;
		instrument1:make_model = "SBE-37" ;
		instrument1:serial_number = "1859723" ;
		instrument1:calibration_date = "2016-03-25" ;
		instrument1:accuracy = "" ;
		instrument1:precision = "" ;
		instrument1:comment = "serial number and calibration dates are bogus" ;
	char platform1 ;
		platform1:long_name = "Underwater Slocum Glider RU07" ;
		platform1:ncei_code = "RU07" ;
		platform1:ioos_code = "urn:ioos:station:NCEI:RU07" ;
		platform1:call_sign = "" ;
		platform1:ices_code = "" ;
		platform1:imo_code = "" ;
		platform1:wmo_code = "4801537" ;
		platform1:comment = "Data is not actually collected from this platform, this is an example." ;
	double crs ;
		crs:grid_mapping_name = "latitude_longitude" ;
		crs:longitude_of_prime_meridian = 0. ;
		crs:semi_major_axis = 6378137. ;
		crs:inverse_flattening = 298.257223563 ;
		crs:epsg_code = "EPSG:4326" ;

// global attributes:
		:instrument = "In Situ/Laboratory Instruments > Profilers/Sounders > > > CTD" ;
		:platform = "In Situ Ocean-based Platforms > > SEAGLIDER" ;
		:title = "Oceanographic and surface meteorological data collected from the Underwater Slocum Glider RU07 by the National Centers for Environmental Information (NCEI) in the Cordell Bank National Marine Sanctuary from 2015-03-25 to 2015-03-25" ;
		:ncei_template_version = "NCEI_NetCDF_TrajectoryProfile_Orthogonal_Template_v2.0" ;
		:Conventions = "CF-1.6, ACDD-1.3" ;
		:naming_authority = "gov.noaa.ncei" ;
		:geospatial_bounds = "LINESTRING (-123.982609294 37.0728913284, -124.22393993 37.5322779699, -124.365223371 38.0392701242, -123.649197851 37.138136132, -123.647583716 37.9526057811, -124.456054314 37.573879111, -123.520624033 37.4778548932, -124.280033663 37.3704533063, -123.770691959 37.2367242254, -124.252704493 37.9785987597)" ;
		:geospatial_bounds_crs = "EPSG:4326" ;
		:geospatial_bounds_vertical_crs = "EPSG:5829" ;
		:creator_type = "person" ;
		:creator_institution = "NCEI" ;
		:publisher_type = "position" ;
		:publisher_institution = "NCEI" ;
		:program = "NCEI-IOOS Data Pipeline" ;
		:date_metadata_modified = "2016-09-22T18:16:16.896731Z" ;
		:product_version = "v1" ;
		:instrument_vocabulary = "GCMD Earth Science Keywords. Version 5.3.3" ;
		:platform_vocabulary = "GCMD Earth Science Keywords. Version 5.3.3" ;
		:summary = "This is an example of the Oceanographic and surface meteorological data collected from the Underwater Slocum Glider RU07 by the National Centers for Environmental Information (NCEI) in the Cordell Bank National Marine Sanctuary from 2015-03-25 to 2015-03-25. The data contained within this file are completely bogus and are generated using the python module numpy.random.rand() function. This file can be used for testing with various applications. The uuid was generated using the uuid python module, invoking the command uuid.uuid4()." ;
		:source = "Python script generate_NCEI_netCDF_template.py with options: {\'template_version\': \'2.0\', \'feature_type\': \'trajectoryProfile\'}" ;
		:featureType = "trajectoryProfile" ;
		:cdm_data_type = "Trajectory" ;
		:standard_name_vocabulary = "CF Standard Name Table v30" ;
		:uuid = "b792c055-1d4e-4bf2-aa68-cdca1826ee1f" ;
		:sea_name = "Cordell Bank National Marine Sanctuary, North Pacific Ocean" ;
		:id = "NCEI_trajectoryProfile_template_v2.0_2016-09-22_181616.896731.nc" ;
		:time_coverage_start = "2015-03-25T22:20:18Z" ;
		:time_coverage_end = "2015-03-25T22:21:48Z" ;
		:time_coverage_resolution = "PT10.S" ;
		:geospatial_lat_min = 37.0728913284183 ;
		:geospatial_lat_max = 38.0392701241658 ;
		:geospatial_lat_units = "degrees_north" ;
		:geospatial_lat_resolution = 0.100634159031136 ;
		:geospatial_lon_min = -124.456054313988 ;
		:geospatial_lon_max = -123.52062403339 ;
		:geospatial_lon_units = "degrees_east" ;
		:geospatial_lon_resolution = -0.030010577643351 ;
		:geospatial_vertical_min = 1 ;
		:geospatial_vertical_max = 4 ;
		:geospatial_vertical_units = "m" ;
		:geospatial_vertical_resolution = 1. ;
		:geospatial_vertical_positive = "down" ;
		:institution = "NCEI" ;
		:creator_name = "Mathew Biddle" ;
		:creator_url = "http://www.nodc.noaa.gov/" ;
		:creator_email = "Mathew.Biddle@noaa.gov" ;
		:project = "NCEI NetCDF templates" ;
		:processing_level = "BOGUS DATA" ;
		:metadata_link = "https://www.nodc.noaa.gov/data/formats/netcdf/v2.0/" ;
		:references = "https://www.nodc.noaa.gov/data/formats/netcdf/v2.0/" ;
		:keywords_vocabulary = "GCMD Earth Science Keywords. Version 5.3.3" ;
		:keywords = "Oceans > Ocean Temperature > Water Temperature, Oceans > Salinity/Density > Salinity" ;
		:acknowledgement = "thanks to the NCEI netCDF working group" ;
		:comment = "This data file is just an example, the data are completely BOGUS!" ;
		:contributor_name = "NCEI" ;
		:contributor_role = "Data Center" ;
		:date_created = "2016-09-22T18:16:16.896731Z" ;
		:date_modified = "2016-09-22T18:16:16.896731Z" ;
		:date_issued = "2016-09-22T18:16:16.896731Z" ;
		:publisher_name = "NCEI Data Manager" ;
		:publisher_email = "ncei.ioos@noaa.gov" ;
		:publisher_url = "http://www.ncei.noaa.gov/" ;
		:license = "Freely available" ;
		:time_coverage_duration = "PT1M30S" ;
		:history = "Tue Sep 27 16:40:22 2016: ncatted -a time_coverage_duration,global,m,c,PT1M30S ./NCEI_trajectoryProfile_template_v2.0_2016-09-22_181616.896731.nc\n",
			"This file was created on 2016-09-22T18:16:16.896731Z" ;
}

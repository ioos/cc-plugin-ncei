netcdf NODC_trajectory_template_v1.1_2016-06-14_125322.975680 {
dimensions:
	maxStrlen64 = 64 ;
	obs = 10 ;
	trajectory = 1 ;
variables:
	int trajectory(trajectory) ;
		trajectory:long_name = "Leg 1 of cruise AVH2016" ;
		trajectory:cf_role = "trajectory_id" ;
		trajectory:_Netcdf4Dimid = 1 ;
	double time(trajectory, obs) ;
		time:_FillValue = -9999. ;
		time:_Netcdf4Dimid = 1 ;
		time:long_name = "Time" ;
		time:standard_name = "time" ;
		time:units = "seconds since 1970-01-01 00:00:00 UTC" ;
		time:axis = "T" ;
		time:calendar = "julian" ;
		time:comment = "This data is BOGUS!!!!!" ;
	double lat(trajectory, obs) ;
		lat:_FillValue = -9999. ;
		lat:_Netcdf4Dimid = 1 ;
		lat:long_name = "Latitude" ;
		lat:standard_name = "latitude" ;
		lat:units = "degrees_north" ;
		lat:axis = "Y" ;
		lat:valid_min = -90. ;
		lat:valid_max = 90. ;
		lat:comment = "This data is BOGUS!!!!!" ;
	double lon(trajectory, obs) ;
		lon:_FillValue = -9999. ;
		lon:_Netcdf4Dimid = 1 ;
		lon:long_name = "Longitude" ;
		lon:standard_name = "longitude" ;
		lon:units = "degrees_east" ;
		lon:axis = "X" ;
		lon:valid_min = -180. ;
		lon:valid_max = 180. ;
		lon:comment = "This data is BOGUS!!!!!" ;
	double z(trajectory, obs) ;
		z:_FillValue = -9999. ;
		z:_Netcdf4Dimid = 1 ;
		z:long_name = "depth of sensor" ;
		z:standard_name = "depth" ;
		z:units = "m" ;
		z:axis = "Z" ;
		z:valid_min = 0. ;
		z:valid_max = 10971. ;
		z:positive = "down" ;
		z:comment = "This data is BOGUS!!!!!" ;
	double sal(trajectory, obs) ;
		sal:_FillValue = -9999. ;
		sal:_Netcdf4Dimid = 1 ;
		sal:long_name = "Salinity" ;
		sal:standard_name = "sea_water_salinity" ;
		sal:nodc_name = "SALINITY" ;
		sal:units = "0.001" ;
		sal:scale_factor = 1. ;
		sal:add_offset = 0. ;
		sal:valid_min = 0. ;
		sal:valid_max = 100. ;
		sal:data_min = 33.0367581975989 ;
		sal:data_max = 33.9316903450518 ;
		sal:coordinates = "time lat lon z" ;
		sal:grid_mapping = "crs" ;
		sal:source = "This data is completely false data, the number was randomly selected" ;
		sal:references = "http://www.numpy.org/" ;
		sal:cell_methods = "time: point longitude: point latitude: point" ;
		sal:platform = "platform1" ;
		sal:instrument = "instrument1" ;
		sal:comment = "This data is BOGUS!!!!!" ;
	double temp(trajectory, obs) ;
		temp:_FillValue = -9999. ;
		temp:long_name = "Temperature" ;
		temp:standard_name = "sea_water_temperature" ;
		temp:nodc_name = "WATER TEMPERATURE" ;
		temp:units = "degree_Celsius" ;
		temp:scale_factor = 1. ;
		temp:add_offset = 0. ;
		temp:valid_min = 0. ;
		temp:valid_max = 100. ;
		temp:data_min = 13.2202028578429 ;
		temp:data_max = 13.8343090768195 ;
		temp:coordinates = "time lat lon z" ;
		temp:grid_mapping = "crs" ;
		temp:source = "This data is completely false data, the number was randomly selected" ;
		temp:references = "http://www.numpy.org/" ;
		temp:cell_methods = "time: point longitude: point latitude: point" ;
		temp:platform = "platform1" ;
		temp:instrument = "instrument1" ;
		temp:comment = "This data is BOGUS!!!!!" ;
	char instrument1(maxStrlen64) ;
		instrument1:comment = "serial number and calibration dates are bogus" ;
		instrument1:calibration_date = "2016-03-25" ;
		instrument1:serial_number = "1859723" ;
		instrument1:long_name = "Seabird SBE 45 MicroTSG Thermosalinograph" ;
		instrument1:nodc_name = "Thermosalinographs" ;
		instrument1:make_model = "SBE-45" ;
	char platform1(maxStrlen64) ;
		platform1:long_name = "Alexander Von Humboldt" ;
		platform1:nodc_code = "ALEXANDER VON HUMBOLDT" ;
		platform1:ioos_code = "urn:ioos:station:NCEI:AlexanderVonHumboldt" ;
		platform1:call_sign = "DFAW" ;
		platform1:imo_code = "8626886" ;
		platform1:comment = "Data is not actually collected from this platform, this is an example." ;
	double crs ;
		crs:grid_mapping_name = "latitude_longitude" ;
		crs:longitude_of_prime_meridian = 0. ;
		crs:semi_major_axis = 6378137. ;
		crs:inverse_flattening = 298.257223563 ;
		crs:epsg_code = "EPSG:4326" ;

// global attributes:
		:instrument = "instrument1" ;
		:platform = "platform1" ;
		:title = "Oceanographic and surface meteorological data collected from the Alexander Von Humboldt by the National Centers for Environmental Information (NCEI) in the Cordell Bank National Marine Sanctuary from 2015-03-25 to 2015-03-25" ;
		:nodc_template_version = "NODC_NetCDF_trajectory_Template_v1.1" ;
		:Conventions = "CF-1.6" ;
		:naming_authority = "gov.noaa.nodc" ;
		:Metadata_Conventions = "Unidata Dataset Discovery v1.0" ;
		:summary = "This is an example of the Oceanographic and surface meteorological data collected from the Alexander Von Humboldt by the National Centers for Environmental Information (NCEI) in the Cordell Bank National Marine Sanctuary from 2015-03-25 to 2015-03-25. The data contained within this file is completely bogus and is generated using the python module numpy.random.rand() function. This file can be used for testing with various applications. The uuid was generated using the uuid python module, invoking the command uuid.uuid4()." ;
		:source = "Python script generate_NCEI_netCDF_template.py with options: {\'template_version\': \'1.1\', \'feature_type\': \'trajectory\'}" ;
		:featureType = "trajectory" ;
		:cdm_data_type = "Trajectory" ;
		:standard_name_vocabulary = "CF Standard Name Table v30" ;
		:uuid = "39eeb570-02cf-4e47-8c8e-f179c68dba61" ;
		:sea_name = "Cordell Bank National Marine Sanctuary, North Pacific Ocean" ;
		:id = "NODC_trajectory_template_v1.1_2016-06-14_125322.975680.nc" ;
		:time_coverage_start = "2015-03-25T22:20:18Z" ;
		:time_coverage_end = "2015-03-25T22:21:48Z" ;
		:time_coverage_resolution = "PT10.S" ;
		:time_coverage_duration = "PT1M30.S" ;
		:geospatial_lat_min = 37.0740875783237 ;
		:geospatial_lat_max = 37.8582057565534 ;
		:geospatial_lat_units = "degrees_north" ;
		:geospatial_lat_resolution = 0.0275870832656982 ;
		:geospatial_lon_min = -124.366980471248 ;
		:geospatial_lon_max = -123.486487373993 ;
		:geospatial_lon_units = "degrees_east" ;
		:geospatial_lon_resolution = 0.076130332683669 ;
		:geospatial_vertical_min = 1.5 ;
		:geospatial_vertical_max = 1.5 ;
		:geospatial_vertical_units = "m" ;
		:geospatial_vertical_resolution = 0. ;
		:geospatial_vertical_positive = "down" ;
		:institution = "NCEI" ;
		:creator_name = "Mathew Biddle" ;
		:creator_url = "http://www.nodc.noaa.gov/" ;
		:creator_email = "Mathew.Biddle@noaa.gov" ;
		:project = "NCEI NetCDF templates" ;
		:processing_level = "BOGUS DATA" ;
		:metadata_link = "https://www.nodc.noaa.gov/data/formats/netcdf/v2.0/" ;
		:keywords_vocabulary = "GCMD Earth Science Keywords. Version 5.3.3" ;
		:keywords = "Oceans > Ocean Temperature > Water Temperature, Oceans > Salinity/Density > Salinity" ;
		:acknowledgement = "thanks to the NCEI netCDF working group" ;
		:comment = "This data file is just an example, the data is completely BOGUS!" ;
		:contributor_name = "NCEI" ;
		:contributor_role = "Data Center" ;
		:date_created = "2016-06-14T12:53:22.975680Z" ;
		:date_modified = "2016-06-14T12:53:22.975680Z" ;
		:date_issued = "2016-06-14T12:53:22.975680Z" ;
		:publisher_name = "NCEI Data Manager" ;
		:publisher_email = "ncei.ioos@noaa.gov" ;
		:publisher_url = "http://www.ncei.noaa.gov/" ;
		:history = "This file was created on 2016-06-14T12:53:22.975680Z" ;
		:license = "Freely available" ;
		:references = "https://www.nodc.noaa.gov/data/formats/netcdf/v2.0/" ;
		:DODS.strlen = 0 ;
}

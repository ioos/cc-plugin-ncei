netcdf BodegaMarineLabBuoyCombined {
dimensions:
	obs = 63242 ;
	timeSeries = 2 ;
variables:
	double time(timeSeries, obs) ;
		time:standard_name = "time" ;
		time:long_name = "Time" ;
		time:units = "seconds since 1970-01-01 00:00:00 UTC" ;
		time:_FillValue = -99999. ;
		time:ancillary_variables = "" ;
		time:comment = "" ;
		time:ioos_category = "Time" ;
		time:calendar = "standard" ;
                time:axis = "T" ;
	float lat(timeSeries) ;
		lat:long_name = "latitude in decimal degrees north" ;
		lat:standard_name = "latitude" ;
		lat:units = "degrees_north" ;
		lat:valid_min = -180. ;
		lat:valid_max = 180. ;
		lat:data_min = 38.0488 ;
		lat:data_max = 38.0488 ;
		lat:instrument = "instrument1" ;
		lat:ancillary_variables = "" ;
		lat:comment = "" ;
		lat:ioos_category = "Location" ;
                lat:axis = "Y" ;
                lat:_FillValue = 0.0f ;
	float lon(timeSeries) ;
		lon:long_name = "longitude in decimal degrees east" ;
		lon:standard_name = "longitude" ;
		lon:units = "degrees_east" ;
		lon:valid_min = -180. ;
		lon:valid_max = 180. ;
		lon:data_min = -123.458 ;
		lon:data_max = -123.458 ;
		lon:instrument = "instrument1" ;
		lon:ancillary_variables = "" ;
		lon:comment = "" ;
		lon:ioos_category = "Location" ;
                lon:axis = "X" ;
                lon:_FillValue = 0.0f ;
	double alt(timeSeries) ;
		alt:long_name = "Height above mean sea level" ;
		alt:standard_name = "altitude" ;
		alt:units = "m" ;
		alt:positive = "up" ;
		alt:valid_min = -10. ;
		alt:valid_max = 0. ;
		alt:data_min = -1.5 ;
		alt:data_max = -1.5 ;
		alt:ancillary_variables = "" ;
		alt:comment = "" ;
		alt:ioos_category = "Location" ;
	     alt:axis = "Z" ;
          alt:_FillValue = 0.0 ;
	int timeSeries(timeSeries) ;
		timeSeries:long_name = "Cordell Bank National Marine Sanctuary (CBNMS) Bodega Marine Lab (BML) Buoy" ;
		timeSeries:cf_role = "timeseries_id" ;
	double temperature(timeSeries, obs) ;
		temperature:long_name = "Water temperature, IPTS-90" ;
		temperature:standard_name = "sea_water_temperature" ;
		temperature:nodc_name = "TEMPERATURE" ;
		temperature:units = "degree_Celsius" ;
		temperature:scale_factor = 1. ;
		temperature:add_offset = 0. ;
		temperature:_FillValue = -99999. ;
		temperature:data_min = 9.8552 ;
		temperature:data_max = 15.8311 ;
		temperature:instrument = "instrument2" ;
		temperature:coordinates = "time lat lon alt" ;
		temperature:source = " " ;
		temperature:references = " " ;
		temperature:ioos_category = "Temperature" ;
		temperature:grid_mapping = "crs" ;
		temperature:ancillary_variables = "temperature_qc" ;
	double salinity(timeSeries, obs) ;
		salinity:long_name = "Salinity, IPSS-78" ;
		salinity:standard_name = "sea_water_salinity" ;
		salinity:nodc_name = "SALINITY" ;
		salinity:units = "0.001" ;
		salinity:scale_factor = 1. ;
		salinity:add_offset = 0. ;
		salinity:_FillValue = -99999. ;
		salinity:data_min = 33.0771 ;
		salinity:data_max = 33.9761 ;
		salinity:instrument = "instrument2" ;
		salinity:coordinates = "time lat lon alt" ;
		salinity:source = " " ;
		salinity:references = " " ;
		salinity:ioos_category = "Salinity" ;
		salinity:grid_mapping = "crs" ;
		salinity:ancillary_variables = "salinity_qc" ;
	double density(timeSeries, obs) ;
		density:long_name = "Density" ;
		density:standard_name = "sea_water_density" ;
		density:nodc_name = "DENSITY" ;
		density:units = "kg m-3" ;
		density:scale_factor = 1. ;
		density:add_offset = 0. ;
		density:_FillValue = -99999. ;
		density:data_min = 24.4722 ;
		density:data_max = 26.1079 ;
		density:instrument = "instrument2" ;
		density:coordinates = "time lat lon alt" ;
		density:source = " " ;
		density:references = " " ;
		density:ioos_category = "Salinity" ;
		density:grid_mapping = "crs" ;
		density:ancillary_variables = "density_qc" ;
	double conductivity(timeSeries, obs) ;
		conductivity:long_name = "Conductivity" ;
		conductivity:standard_name = "sea_water_electrical_conductivity" ;
		conductivity:nodc_name = "CONDUCTIVITY" ;
		conductivity:units = "S m-1" ;
		conductivity:scale_factor = 1. ;
		conductivity:add_offset = 0. ;
		conductivity:_FillValue = -99999. ;
		conductivity:data_min = 3.6799 ;
		conductivity:data_max = 4.18236 ;
		conductivity:instrument = "instrument2" ;
		conductivity:coordinates = "time lat lon alt" ;
		conductivity:source = " " ;
		conductivity:references = " " ;
		conductivity:ioos_category = "Salinity" ;
		conductivity:grid_mapping = "crs" ;
		conductivity:ancillary_variables = "conductivity_qc" ;
	double turbidity(timeSeries, obs) ;
		turbidity:long_name = "Raw Turbidity" ;
		turbidity:nodc_name = "TURBIDITY" ;
		turbidity:units = "NTU" ;
		turbidity:scale_factor = 1. ;
		turbidity:add_offset = 0. ;
		turbidity:_FillValue = -99999. ;
		turbidity:valid_min = 0. ;
		turbidity:valid_max = 4200. ;
		turbidity:data_min = 71. ;
		turbidity:data_max = 2013. ;
		turbidity:instrument = "instrument3" ;
		turbidity:coordinates = "time lat lon alt" ;
		turbidity:source = " " ;
		turbidity:references = " " ;
		turbidity:grid_mapping = "crs" ;
		turbidity:ancillary_variables = "turbidity_qc" ;
		turbidity:ioos_category = "Optical Properties" ;
		turbidity:comment = "Nephelometric Turbidity Unit (NTU) -specs as reported by Wetlabs for concentration; factory calibration scale factor is 0.0060 (NTU soln value was 2189 counts, cal temp 21.5 deg C), dark counts - 45 counts, max output - 4121 counts, resolution, 0.7 counts, for conversion to concentration if desired. Last factory cal for this period: 6/30/2006 (ECO SN 524)." ;
	double fluorescence(timeSeries, obs) ;
		fluorescence:long_name = "Raw Fluorescence" ;
		fluorescence:nodc_name = "FLUORESCENCE" ;
		fluorescence:units = "1" ;
		fluorescence:scale_factor = 1. ;
		fluorescence:add_offset = 0. ;
		fluorescence:_FillValue = -99999. ;
		fluorescence:valid_min = 0. ;
		fluorescence:valid_max = 4200. ;
		fluorescence:data_min = 104. ;
		fluorescence:data_max = 1761. ;
		fluorescence:instrument = "instrument3" ;
		fluorescence:coordinates = "time lat lon alt" ;
		fluorescence:source = " " ;
		fluorescence:references = " " ;
		fluorescence:grid_mapping = "crs" ;
		fluorescence:ancillary_variables = "fluorescence_qc" ;
		fluorescence:ioos_category = "Ocean Color " ;
	int platform1 ;
		platform1:long_name = "Station 46095. Cordell Bank Buoy" ;
		platform1:nodc_name = "FIXED PLATFORM, MOORINGS" ;
		platform1:call_sign = "" ;
		platform1:ices_code = "" ;
		platform1:imo_code = "" ;
		platform1:wmo_code = "46095" ;
		platform1:comment = "" ;
	int temperature_qc(timeSeries, obs) ;
		temperature_qc:standard_name = "sea_water_temperature status_flag" ;
		temperature_qc:long_name = "Temperature QC Flag" ;
		temperature_qc:flag_values = 0, 1, 2, 9 ;
		temperature_qc:flag_meanings = "no_known_bad_data known_bad_data suspicous_data missing_data" ;
		temperature_qc:_FillValue = -99999 ;
		temperature_qc:data_min = 0. ;
		temperature_qc:data_max = 1. ;
		temperature_qc:valid_range = 0., 9. ;
		temperature_qc:coordinates = "time lat lon alt" ;
		temperature_qc:comment = "" ;
	int salinity_qc(timeSeries, obs) ;
		salinity_qc:standard_name = "sea_water_salinity status_flag" ;
		salinity_qc:long_name = "Salinity QC Flag" ;
		salinity_qc:flag_values = 0, 1, 2, 9 ;
		salinity_qc:flag_meanings = "no_known_bad_data known_bad_data suspicous_data missing_data" ;
		salinity_qc:_FillValue = -99999 ;
		salinity_qc:data_min = 0. ;
		salinity_qc:data_max = 0. ;
		salinity_qc:valid_range = 0., 9. ;
		salinity_qc:coordinates = "time lat lon alt" ;
		salinity_qc:comment = "" ;
	int density_qc(timeSeries, obs) ;
		density_qc:standard_name = "sea_water_density status_flag" ;
		density_qc:long_name = "Density QC Flag" ;
		density_qc:flag_values = 0, 1, 2, 9 ;
		density_qc:flag_meanings = "no_known_bad_data known_bad_data suspicous_data missing_data" ;
		density_qc:_FillValue = -99999 ;
		density_qc:data_min = 0. ;
		density_qc:data_max = 0. ;
		density_qc:valid_range = 0., 9. ;
		density_qc:coordinates = "time lat lon alt" ;
		density_qc:comment = "" ;
	int conductivity_qc(timeSeries, obs) ;
		conductivity_qc:standard_name = "sea_water_electrical_conductivity status_flag" ;
		conductivity_qc:long_name = "Conductivity QC Flag" ;
		conductivity_qc:flag_values = 0, 1, 2, 9 ;
		conductivity_qc:flag_meanings = "no_known_bad_data known_bad_data suspicous_data missing_data" ;
		conductivity_qc:_FillValue = -99999 ;
		conductivity_qc:data_min = 0. ;
		conductivity_qc:data_max = 0. ;
		conductivity_qc:valid_range = 0., 9. ;
		conductivity_qc:coordinates = "time lat lon alt" ;
		conductivity_qc:comment = "" ;
	int turbidity_qc(timeSeries, obs) ;
		turbidity_qc:long_name = "Raw Turbidity QC Flag" ;
		turbidity_qc:flag_values = 0, 1, 2, 9 ;
		turbidity_qc:flag_meanings = "no_known_bad_data known_bad_data suspicous_data missing_data" ;
		turbidity_qc:_FillValue = -99999 ;
		turbidity_qc:data_min = 0. ;
		turbidity_qc:data_max = 2. ;
		turbidity_qc:valid_range = 0., 9. ;
		turbidity_qc:coordinates = "time lat lon alt" ;
		turbidity_qc:comment = "" ;
	int fluorescence_qc(timeSeries, obs) ;
		fluorescence_qc:long_name = "Raw Fluorescence QC Flag" ;
		fluorescence_qc:flag_values = 0, 1, 2, 9 ;
		fluorescence_qc:flag_meanings = "no_known_bad_data known_bad_data suspicous_data missing_data" ;
		fluorescence_qc:_FillValue = -99999 ;
		fluorescence_qc:data_min = 0. ;
		fluorescence_qc:data_max = 2. ;
		fluorescence_qc:valid_range = 0., 9. ;
		fluorescence_qc:coordinates = "time lat lon alt" ;
		fluorescence_qc:comment = "" ;
	int instrument1(timeSeries) ;
		instrument1:long_name = "Worldwide GPS Satellite Tracker" ;
		instrument1:nodc_name = "GPS" ;
		instrument1:make_model = "SX1" ;
		instrument1:serial_number = "" ;
		instrument1:calibration_date = "" ;
		instrument1:comment = "" ;
	int instrument2(timeSeries) ;
		instrument2:long_name = "Seabird 37 Microcat" ;
		instrument2:nodc_name = "CTD" ;
		instrument2:make_model = "SBE-37" ;
		instrument2:serial_number = "" ;
		instrument2:calibration_date = "" ;
		instrument2:comment = "" ;
	int instrument3(timeSeries) ;
		instrument3:long_name = "Wetlabs ECO Fluorescence and Turbidity Sensor (ECO-FLNTUSB)" ;
		instrument3:nodc_name = "fluorometer, Turbidity Meter" ;
		instrument3:make_model = "FLNTUSB" ;
		instrument3:scale_factor_fl = 0.0121 ;
		instrument3:dark_counts_fl = 44. ;
		instrument3:max_output_fl = 4121. ;
		instrument3:resolution_fl = "0.8 counts" ;
		instrument3:scale_factor_tu = 0.006 ;
		instrument3:dark_counts_tu = 45. ;
		instrument3:NTU_solution_value = 2189. ;
		instrument3:max_output_tu = 4121. ;
		instrument3:resolution_tu = "0.7 counts" ;
		instrument3:cal_temp = "21.5 degC" ;
		instrument3:comment = "" ;
		instrument3:serial_number = 524. ;
		instrument3:calibration_date = "06/30/2006" ;
	double ht_wgs84(timeSeries) ;
		ht_wgs84:long_name = "Height above WGS 84" ;
		ht_wgs84:standard_name = "height_above_reference_ellipsoid" ;
		ht_wgs84:units = "m" ;
		ht_wgs84:data_min = -34.023998260498 ;
		ht_wgs84:data_max = -34.023998260498 ;
		ht_wgs84:ioos_category = "" ;
		ht_wgs84:ellipsoid_name = "WGS 84" ;
		ht_wgs84:_FillValue = -99999. ;
		ht_wgs84:comment = "" ;
	double ht_mllw(timeSeries) ;
		ht_mllw:long_name = "Height above mean lower low water" ;
		ht_mllw:standard_name = "water_surface_height_above_reference_datum" ;
		ht_mllw:data_min = -0.549000024795532 ;
		ht_mllw:data_max = -0.549000024795532 ;
		ht_mllw:ioos_category = "" ;
		ht_mllw:water_surface_reference_datum_altitude = "lower low water datum" ;
		ht_mllw:_FillValue = -99999. ;
		ht_mllw:comment = "Mean Lower Low Water - The average of the lower low water height of each tidal day observed over the National Tidal Datum Epoch. As defined by NOAA Tides and Currents (http://tidesandcurrents.noaa.gov/datum_options.html)" ;
	int crs ;
		crs:grid_mapping_name = "latitude_longitude" ;
		crs:longitude_of_prime_meridian = 0. ;
		crs:semi_major_axis = 6378137. ;
		crs:inverse_flattening = 298.257223563 ;
		crs:epsg_code = "EPSG:4326" ;

// global attributes:
		:title = "Data collected from Cordell Bank, California, USA, by CBNMS and BML" ;
		:summary = "These seawater data are collected by a moored fluorescence and turbidity instrument operated at Cordell Bank, California, USA, by CBNMS and BML. Beginning on 2008-04-23, fluorescence and turbidity measurements were collected using a Wetlabs ECO Fluorescence and Turbidity Sensor (ECO-FLNTUSB). The instrument depth of the water quality sensors was 01.0 meter, in an overall water depth of 85 meters (both relative to Mean Sea Level, MSL). The measurements reflect a 10 minute sampling interval." ;
		:summary2 = "These seawater data are collected by a moored fluorescence and turbidity instrument operated at Cordell Bank, California, USA, by CBNMS and BML. Beginning on 2008-04-23, fluorescence and turbidity measurements were collected using a Wetlabs ECO Fluorescence and Turbidity Sensor (ECO-FLNTUSB). The instrument depth of the water quality sensors was 01.0 meter, in an overall water depth of 85 meters (both relative to Mean Sea Level, MSL). The measurements reflect a 10 minute sampling interval." ;
		:id = "CBNMS_BML_Bouy_CTD_SFX_combined_v2" ;
		:uuid = "ab0cc5bf-488d-4a65-87d2-90e6471ab21f" ;
		:naming_authority = "gov.noaa.nodc" ;
		:time_coverage_start1 = "2008-07-28 17:30:00 UTC" ;
		:time_coverage_end1 = "2008-09-10 15:31:00 UTC" ;
		:time_coverage_start2 = "2008-07-28 17:33:05 UTC" ;
		:time_coverage_end2 = "2008-09-10 16:33:05 UTC" ;
		:time_coverage_resolution1 = "P1M12DT22H1M" ;
		:time_coverage_resolution2 = "P1M12DT23H" ;
		:platform = "platform1" ;
		:geospatial_lon_max = -123.458000183105 ;
		:geospatial_lon_min = -123.458000183105 ;
		:geospatial_lon_units = "degree_east" ;
		:geospatial_lon_resolution = "point" ;
		:geospatial_lat_max = 38.0488014221191 ;
		:geospatial_lat_min = 38.0488014221191 ;
		:geospatial_lat_units = "degree_north" ;
		:geospatial_lat_resolution = "point" ;
		:geospatial_vertical_min = -1.5 ;
		:geospatial_vertical_max = -1.5 ;
		:geospatial_vertical_positive = "up" ;
		:geospatial_vertical_units = "m" ;
		:geospatial_vertical_reference = "mean_sea_level" ;
		:area = "Cordell Bank National Marine Sanctuary, CA, USA" ;
		:creator_name = "Data Manager (bmldata@ucdavis.edu)" ;
		:infoURL = "http://portal.ncddc.noaa.gov" ;
		:institution = "National Marine Sanctuary Program (NMS), Cordell Bank National Marine Sanctuary (CBNMS) and Bodega Marine Laboratory, University of California Davis" ;
		:institution_url = "http://bml.ucdavis.edu" ;
		:institution_dods_url = "http://bml.ucdavis.edu" ;
		:creator_email = "Data Manager (bmldata@ucdavis.edu)" ;
		:creator_url = "http://bml.ucdavis.edu" ;
		:project = "CBNMS" ;
		:source = "moored platform observation - fixed altitude" ;
		:acknowledgment = "" ;
		:processing_level = "Quality Controlled" ;
		:keywords = "EARTH SCIENCE > Oceans > Ocean Pressure > Water Pressure, EARTH SCIENCE > Oceans > Salinity/Density > Density, EARTH SCIENCE > Oceans > Ocean Temperature > Water Temperature, EARTH SCIENCE > Oceans > Salinity/Density > Conductivity, EARTH SCIENCE > Oceans > Salinity/Density > Salinity" ;
		:keywords_vocabulary = "GCMD Earth Science Keywords. Version 5.3.3" ;
		:standard_name_vocabulary = "NetCDF Climate and Forecast (CF) Metadata Convention Standard Name Table v23" ;
		:comment = "" ;
		:contributor_name = "Megan Sheridan" ;
		:contributor_role = "Staff Research Associate at UC Davis/Bodega Marine Lab" ;
		:originator_files = "NMS_CBM_SFX_2008.nc and NMS_CBM_CTD_2008.nc" ;
		:cdm_data_type = "Station" ;
		:date_created = "24-Apr-2012" ;
		:date_modified = "24-Apr-2012" ;
		:publisher_name = "US NATIONAL OCEANOGRAPHIC DATA CENTER " ;
		:publisher_url = "http://www.nodc.noaa.gov/" ;
		:publisher_email = "NODC.Services@noaa.gov" ;
		:featureType = "timeSeries" ;
		:history = "2011-03-17 23:17:49 UTC: File created at 2011-03-17 23:17:49 UTC edited on 24-Apr-2012 Time units updated on 01-Jan-2013, time units were incorrectly listed as hours since 1970-01-01 00:00:00 UTC instead of seconds since 1970-01-01 00:00:00 UTC; dimensions for station_name were incorrect and have been adjusted to (timeSeries, name_strlen) instead of name_strlen. Conventions gloabal attribute has been adjusted to correctly document the current version of CF used in this example. Values for station_name were adjusted to Cordell_1 and Cordell_2." ;
		:Conventions = "CF-1.6" ;
		:Metadata_Conventions = "Unidata Dataset Discovery v1.0" ;
		:nodc_template_version = "NODC_NetCDF_TimeSeries_Incomplete_Template_v1.1" ;
		:metadata_link = "" ;
}

netcdf BodegaMarineLabBuoy {
dimensions:
	timeSeries = 17 ;
	time = 63242 ;
variables:
	double time(time) ;
		time:standard_name = "time" ;
		time:long_name = "Time" ;
		time:units = "seconds since 1970-01-01 00:00:00 UTC" ;
		time:axis = "T" ;
		time:ancillary_variables = "" ;
		time:comment = "" ;
		time:ioos_category = "Time" ;
		time:calendar = "standard" ;
	float lat ;
		lat:long_name = "latitude in decimal degrees north" ;
		lat:standard_name = "latitude" ;
		lat:units = "degrees_north" ;
		lat:data_min = 38.0488 ;
		lat:data_max = 38.0488 ;
		lat:instrument = "instrument1" ;
		lat:ancillary_variables = "" ;
		lat:comment = "" ;
		lat:ioos_category = "Location" ;
                lat:axis = "Y" ;
                lat:_FillValue = 0.0f ;
                lat:valid_min = -90.0 ;
                lat:valid_max = 90.0 ; 
	float lon ;
		lon:long_name = "longitude in decimal degrees east" ;
		lon:standard_name = "longitude" ;
		lon:units = "degrees_east" ;
		lon:data_min = -123.458 ;
		lon:data_max = -123.458 ;
		lon:instrument = "instrument1" ;
		lon:ancillary_variables = "" ;
		lon:comment = "" ;
		lon:ioos_category = "Location" ;
                lon:axis ="X" ;
                lon:_FillValue = 0.0f ;
                lon:valid_min = -180.0 ;
                lon:valid_max = 180.0 ; 
	double alt ;
		alt:long_name = "Height above mean sea level" ;
		alt:standard_name = "altitude" ;
		alt:units = "m" ;
		alt:positive = "up" ;
		alt:data_min = -1.5 ;
		alt:data_max = -1.5 ;
		alt:ancillary_variables = "" ;
		alt:comment = "" ;
		alt:ioos_category = "Location" ;
                alt:axis = "Z" ;
                alt:_FillValue = 0.0 ;
                alt:valid_min = -200.0 ;
                alt:valid_max = 0.0 ; 
	char timeSeries(timeSeries) ;
		timeSeries:long_name = "Cordell Bank National Marine Sanctuary (CBNMS) Bodega Marine Lab (BML) Buoy" ;
		timeSeries:cf_role = "timeseries_id" ;
	double temperature(time) ;
		temperature:long_name = "Water temperature, IPTS-90" ;
		temperature:standard_name = "sea_water_temperature" ;
		temperature:nodc_name = "TEMPERATURE" ;
		temperature:units = "degree_Celsius" ;
		temperature:scale_factor = 1. ;
		temperature:add_offset = 0. ;
		temperature:_FillValue = -99999. ;
		temperature:data_min = 9.8552 ;
		temperature:data_max = 15.8311 ;
		temperature:instrument = "instrument2" ;
		temperature:coordinates = "time lat lon alt" ;
		temperature:source = " " ;
		temperature:references = " " ;
		temperature:ioos_category = "Temperature" ;
		temperature:grid_mapping = "crs" ;
		temperature:ancillary_variables = "temperature_qc" ;
                temperature:valid_min = -200.0 ;
                temperature:valid_max = 0.0 ;
                temperature:comment = "comment" ;
	double salinity(time) ;
		salinity:long_name = "Salinity, IPSS-78" ;
		salinity:standard_name = "sea_water_salinity" ;
		salinity:nodc_name = "SALINITY" ;
		salinity:units = "0.001" ;
		salinity:scale_factor = 1. ;
		salinity:add_offset = 0. ;
		salinity:_FillValue = -99999. ;
		salinity:data_min = 33.0771 ;
		salinity:data_max = 33.9761 ;
		salinity:instrument = "instrument2" ;
		salinity:coordinates = "time lat lon alt" ;
		salinity:source = " " ;
		salinity:references = " " ;
		salinity:ioos_category = "Salinity" ;
		salinity:grid_mapping = "crs" ;
		salinity:ancillary_variables = "salinity_qc" ;
                salinity:valid_min = -200.0 ;
                salinity:valid_max = 0.0 ; 
                salinity:comment = "comment" ;
	double density(time) ;
		density:long_name = "Density" ;
		density:standard_name = "sea_water_density" ;
		density:nodc_name = "DENSITY" ;
		density:units = "kg m-3" ;
		density:scale_factor = 1. ;
		density:add_offset = 0. ;
		density:_FillValue = -99999. ;
		density:data_min = 24.4722 ;
		density:data_max = 26.1079 ;
		density:instrument = "instrument2" ;
		density:coordinates = "time lat lon alt" ;
		density:source = " " ;
		density:references = " " ;
		density:ioos_category = "Salinity" ;
		density:grid_mapping = "crs" ;
		density:ancillary_variables = "density_qc" ;
                density:valid_min = -200.0 ;
                density:valid_max = 0.0 ; 
                density:comment = "comment" ;
	double conductivity(time) ;
		conductivity:long_name = "Conductivity" ;
		conductivity:standard_name = "sea_water_electrical_conductivity" ;
		conductivity:nodc_name = "CONDUCTIVITY" ;
		conductivity:units = "S m-1" ;
		conductivity:scale_factor = 1. ;
		conductivity:add_offset = 0. ;
		conductivity:_FillValue = -99999. ;
		conductivity:data_min = 3.6799 ;
		conductivity:data_max = 4.18236 ;
		conductivity:instrument = "instrument2" ;
		conductivity:coordinates = "time lat lon alt" ;
		conductivity:source = " " ;
		conductivity:references = " " ;
		conductivity:ioos_category = "Salinity" ;
		conductivity:grid_mapping = "crs" ;
		conductivity:ancillary_variables = "conductivity_qc" ;
                conductivity:valid_min = -200.0 ;
                conductivity:valid_max = 0.0 ; 
                conductivity:comment = "comment" ;
	int platform1 ;
		platform1:long_name = "Station 46095. Cordell Bank Buoy" ;
		platform1:nodc_name = "FIXED PLATFORM, MOORINGS" ;
		platform1:call_sign = "" ;
		platform1:ices_code = "" ;
		platform1:imo_code = "" ;
		platform1:wmo_code = "46095" ;
		platform1:comment = "" ;
        platform1:nodc_code = "" ;
	int temperature_qc(time) ;
		temperature_qc:standard_name = "sea_water_temperature status_flag" ;
		temperature_qc:long_name = "Temperature QC Flag" ;
		temperature_qc:flag_values = 0, 1, 2, 9 ;
		temperature_qc:flag_meanings = "no_known_bad_data, known_bad_data, suspicous_data, missing_data" ;
		temperature_qc:data_min = 0. ;
		temperature_qc:data_max = 1. ;
		temperature_qc:valid_range = 0., 9. ;
		temperature_qc:coordinates = "time lat lon alt" ;
		temperature_qc:_FillValue = 0 ;
		temperature_qc:comment = "" ;
		temperature_qc:references = " " ;
	int salinity_qc(time) ;
		salinity_qc:standard_name = "sea_water_salinity status_flag" ;
		salinity_qc:long_name = "Salinity QC Flag" ;
		salinity_qc:flag_values = 0, 1, 2, 9 ;
		salinity_qc:flag_meanings = "no_known_bad_data, known_bad_data, suspicous_data, missing_data" ;
		salinity_qc:data_min = 0. ;
		salinity_qc:data_max = 0. ;
		salinity_qc:valid_range = 0., 9. ;
		salinity_qc:coordinates = "time lat lon alt" ;
		salinity_qc:_FillValue = 0 ;
		salinity_qc:comment = "" ;
		salinity_qc:references = " " ;
	int density_qc(time) ;
		density_qc:standard_name = "sea_water_density status_flag" ;
		density_qc:long_name = "Density QC Flag" ;
		density_qc:flag_values = 0, 1, 2, 9 ;
		density_qc:flag_meanings = "no_known_bad_data, known_bad_data, suspicous_data, missing_data" ;
		density_qc:data_min = 0. ;
		density_qc:data_max = 0. ;
		density_qc:valid_range = 0., 9. ;
		density_qc:coordinates = "time lat lon alt" ;
		density_qc:_FillValue = 0 ;
		density_qc:comment = "" ;
		density_qc:references = " " ;
	int conductivity_qc(time) ;
		conductivity_qc:standard_name = "sea_water_electrical_conductivity status_flag" ;
		conductivity_qc:long_name = "Conductivity QC Flag" ;
		conductivity_qc:flag_values = 0, 1, 2, 9 ;
		conductivity_qc:flag_meanings = "no_known_bad_data, known_bad_data, suspicous_data, missing_data" ;
		conductivity_qc:data_min = 0. ;
		conductivity_qc:data_max = 0. ;
		conductivity_qc:valid_range = 0., 9. ;
		conductivity_qc:coordinates = "time lat lon alt" ;
		conductivity_qc:_FillValue = 0 ;
		conductivity_qc:comment = "" ;
		conductivity_qc:references = " " ;
	int instrument1 ;
		instrument1:long_name = "Worldwide GPS Satellite Tracker" ;
		instrument1:nodc_name = "GPS" ;
		instrument1:make_model = "SX1" ;
		instrument1:serial_number = "" ;
		instrument1:calibration_date = "" ;
		instrument1:comment = "GPS tracker" ;
	int instrument2 ;
		instrument2:long_name = "Seabird 37 Microcat" ;
		instrument2:nodc_name = "CTD" ;
		instrument2:make_model = "SBE-37" ;
		instrument2:serial_number = "" ;
		instrument2:calibration_date = "" ;
		instrument2:comment = "CTD" ;
	double ht_wgs84 ;
		ht_wgs84:long_name = "Height above WGS 84" ;
		ht_wgs84:standard_name = "height_above_reference_ellipsoid" ;
		ht_wgs84:units = "m" ;
		ht_wgs84:data_min = -34.023998260498 ;
		ht_wgs84:data_max = -34.023998260498 ;
		ht_wgs84:ioos_category = "" ;
		ht_wgs84:ellipsoid_name = "WGS 84" ;
		ht_wgs84:_FillValue = -99999. ;
		ht_wgs84:comment = "" ;
	double ht_mllw ;
		ht_mllw:long_name = "Height above mean lower low water" ;
		ht_mllw:standard_name = "water_surface_height_above_reference_datum" ;
		ht_mllw:data_min = -0.549000024795532 ;
		ht_mllw:data_max = -0.549000024795532 ;
		ht_mllw:ioos_category = "" ;
		ht_mllw:water_surface_reference_datum_altitude = "lower low water datum" ;
		ht_mllw:_FillValue = -99999. ;
		ht_mllw:comment = "Mean Lower Low Water - The average of the lower low water height of each tidal day observed over the National Tidal Datum Epoch. As defined by NOAA Tides and Currents (http://tidesandcurrents.noaa.gov/datum_options.html)" ;
	int crs ;
		crs:grid_mapping_name = "latitude_longitude" ;
		crs:longitude_of_prime_meridian = 0. ;
		crs:semi_major_axis = 6378137. ;
		crs:inverse_flattening = 298.257223563 ;
		crs:epsg_code = "EPSG:4326" ;

// global attributes:
		:title = "Data collected from Cordell Bank, California, USA, by CBNMS and BML" ;
		:summary = "These seawater data are collected by a moored fluorescence and turbidity instrument operated at Cordell Bank, California, USA, by CBNMS and BML. Beginning on 2008-04-23, fluorescence and turbidity measurements were collected using a Wetlabs ECO Fluorescence and Turbidity Sensor (ECO-FLNTUSB). The instrument depth of the water quality sensors was 01.0 meter, in an overall water depth of 85 meters (both relative to Mean Sea Level, MSL). The measurements reflect a 10 minute sampling interval." ;
		:id = "CBNMS_BML_Bouy_CTD_v2" ;
		:uuid = "846348cd-423f-4358-b9c3-e5e1bf92bc40" ;
		:naming_authority = "gov.noaa.nodc" ;
		:time_coverage_start = "2008-07-28T17:30:00Z" ;
		:time_coverage_end = "2008-09-10T15:31:00Z" ;
		:time_coverage_resolution = "P1M12DT22H28M" ;
		:platform = "platform1" ;
		:geospatial_lon_max = -123.458000183105 ;
		:geospatial_lon_min = -123.458000183105 ;
		:geospatial_lon_units = "degrees_east" ;
		:geospatial_lon_resolution = "point" ;
		:geospatial_lat_max = 38.0488014221191 ;
		:geospatial_lat_min = 38.0488014221191 ;
		:geospatial_lat_units = "degrees_north" ;
		:geospatial_lat_resolution = "point" ;
		:geospatial_vertical_min = -1.5 ;
		:geospatial_vertical_max = -1.5 ;
		:geospatial_vertical_positive = "up" ;
		:geospatial_vertical_units = "m" ;
        :geospatial_vertical_resolution = "point" ;
		:geospatial_vertical_reference = "mean_sea_level" ;
		:area = "Cordell Bank National Marine Sanctuary, CA, USA" ;
		:creator_name = "Data Manager (bmldata@ucdavis.edu)" ;
		:infoURL = "http://portal.ncddc.noaa.gov" ;
		:institution = "National Marine Sanctuary Program (NMS), Cordell Bank National Marine Sanctuary (CBNMS) and Bodega Marine Laboratory, University of California Davis" ;
		:institution_url = "http://bml.ucdavis.edu" ;
		:institution_dods_url = "http://bml.ucdavis.edu" ;
		:creator_email = "Data Manager (bmldata@ucdavis.edu)" ;
		:creator_url = "http://bml.ucdavis.edu" ;
		:project = "CBNMS" ;
		:source = "moored platform observation - fixed altitude" ;
		:acknowledgment = "Data collected from Cordell Bank, California, USA, by CBNMS and BML" ;
		:processing_level = "Quality Controlled" ;
		:keywords = "EARTH SCIENCE > Oceans > Ocean Pressure > Water Pressure, EARTH SCIENCE > Oceans > Salinity/Density > Density, EARTH SCIENCE > Oceans > Ocean Temperature > Water Temperature, EARTH SCIENCE > Oceans > Salinity/Density > Conductivity, EARTH SCIENCE > Oceans > Salinity/Density > Salinity" ;
		:keywords_vocabulary = "GCMD Earth Science Keywords. Version 5.3.3" ;
		:standard_name_vocabulary = "NetCDF Climate and Forecast (CF) Metadata Convention Standard Name Table v23" ;
		:comment = "This dataset is used by the compliance checker as a test dataset" ;
		:contributor_name = "Megan Sheridan" ;
		:contributor_role = "Staff Research Associate at UC Davis/Bodega Marine Lab" ;
		:originator_files = "NMS_CBM_CTD_2008.nc" ;
		:cdm_data_type = "Station" ;
		:date_created = "2012-04-24" ;
		:date_modified = "2012-04-24" ;
		:publisher_name = "US NATIONAL OCEANOGRAPHIC DATA CENTER " ;
		:publisher_url = "http://www.nodc.noaa.gov/" ;
		:publisher_email = "NODC.Services@noaa.gov" ;
		:featureType = "timeSeries" ;
		:history = "2011-03-17 23:17:49 UTC: File created at 2011-03-17 23:17:49 UTC edited on 24-Apr-2012 Time units updated on 01-Jan-2013, time units were incorrectly listed as hours since 1970-01-01 00:00:00 UTC instead of seconds since 1970-01-01 00:00:00 UTC" ;
		:Conventions = "CF-1.6" ;
		:Metadata_Conventions = "Unidata Dataset Discovery v1.0" ;
		:nodc_template_version = "NODC_NetCDF_TimeSeries_Orthogonal_Template_v1.1" ;
		:metadata_link = "http://google.com" ;
        :sea_name = "Coastal Waters of California" ;
        :license = "This data is a reference dataset for the IOOS compliance checker for testing purposes ONLY." ;
        :references = "A reference" ; 
}

netcdf aoml_tsg {
dimensions:
	trajectory = 1 ;
	obs = 2880 ;
variables:
	int trajectory(trajectory) ;
		trajectory:long_name = "trajectory name" ;
		trajectory:cf_role = "trajectory_id" ;
	int time(trajectory, obs) ;
		time:long_name = "time" ;
		time:standard_name = "time" ;
		time:units = "seconds since 2008-06-15 00:00:00 0:00" ;
		time:instrument = "GPS" ;
		time:axis = "T" ;
		time:ancillary_variables = "flag_b, flag_e" ;
                time:calendar = "julian" ;
                time:_FillValue = 0.0f ;
	double lat(trajectory, obs) ;
		lat:long_name = "latitude" ;
		lat:standard_name = "latitude" ;
		lat:units = "degrees_north" ;
		lat:valid_min = -90. ;
		lat:valid_max = 90. ;
		lat:instrument = "GPS" ;
		lat:grid_mapping = "crs" ;
		lat:ancillary_variables = "flag_c, flag_d, flag_e" ;
	double lon(trajectory, obs) ;
		lon:long_name = "longitude" ;
		lon:standard_name = "longitude" ;
		lon:units = "degrees_east" ;
		lon:valid_min = -180. ;
		lon:valid_max = 180. ;
		lon:instrument = "GPS" ;
		lon:grid_mapping = "crs" ;
		lon:ancillary_variables = "flag_c, flag_d, flag_e" ;
	double intp(trajectory, obs) ;
		intp:long_name = "internal thermosalinograph temperature" ;
		intp:units = "degree_Celsius" ;
		intp:_FillValue = -99999. ;
		intp:valid_min = -2.5 ;
		intp:valid_max = 45. ;
		intp:instrument = "tsg" ;
		intp:coordinates = "time lat lon" ;
		intp:grid_mapping = "crs" ;
		intp:nodc_name = "temperature" ;
		intp:ancillary_variables = "flag_f, flag_g, flag_h, flag_i, flag_j, flag_k, flag_l" ;
	double sal(trajectory, obs) ;
		sal:long_name = "thermosalinograph salinity" ;
		sal:standard_name = "sea_water_salinity" ;
		sal:units = "1e-3" ;
		sal:_FillValue = -99999. ;
		sal:valid_min = 0. ;
		sal:valid_max = 60. ;
		sal:instrument = "tsg" ;
		sal:coordinates = "time lat lon" ;
		sal:grid_mapping = "crs" ;
		sal:comment = "Data values are reported in PSU." ;
		sal:nodc_name = "salinity" ;
		sal:ancillary_variables = "flag_f, flag_g, flag_h, flag_i, flag_j, flag_k, flag_l" ;
	double cond(trajectory, obs) ;
		cond:long_name = "thermosalinograph conductivity" ;
		cond:standard_name = "sea_water_electrical_conductivity" ;
		cond:units = "S m-1" ;
		cond:_FillValue = -99999. ;
		cond:valid_min = 0. ;
		cond:valid_max = 6. ;
		cond:instrument = "tsg" ;
		cond:coordinates = "time lat lon" ;
		cond:grid_mapping = "crs" ;
		cond:nodc_name = "conductivity" ;
	double ext(trajectory, obs) ;
		ext:long_name = "thermistor water temperature" ;
		ext:standard_name = "sea_water_temperature" ;
		ext:units = "degree_Celsius" ;
		ext:_FillValue = -99999. ;
		ext:valid_min = -2.5 ;
		ext:valid_max = 45. ;
		ext:instrument = "tmsr" ;
		ext:coordinates = "time lat lon" ;
		ext:grid_mapping = "crs" ;
		ext:nodc_name = "temperature" ;
		ext:ancillary_variables = "flag_f, flag_g, flag_h, flag_i, flag_j, flag_k, flag_l" ;
	double sst(trajectory, obs) ;
		sst:long_name = "sea surface temperature" ;
		sst:standard_name = "sea_water_temperature" ;
		sst:units = "degree_Celsius" ;
		sst:_FillValue = -99999. ;
		sst:valid_min = -2.5 ;
		sst:valid_max = 45. ;
		sst:instrument = "sstr" ;
		sst:coordinates = "time lat lon" ;
		sst:grid_mapping = "crs" ;
		sst:nodc_name = "sea surface temperature" ;
		sst:ancillary_variables = "flag_f, flag_g, flag_h, flag_i, flag_j, flag_k, flag_l" ;
	byte plt(trajectory) ;
		plt:long_name = "David Starr Jordan" ;
		plt:call_sign = "WTDK" ;
		plt:imo_code = "7333195" ;
		plt:platform_technician_email_address = "ChiefET.Jordan@noaa.gov" ;
		plt:platform_technician_alternate_email_address = "n/a" ;
		plt:ancillary_variables = "flag_a" ;
	byte tsg(trajectory) ;
		tsg:long_name = "underway thermosalinograph" ;
		tsg:nodc_name = "thermosalinographs" ;
		tsg:make_model = "SBE-21" ;
		tsg:serial_number = "2118494-2647" ;
		tsg:calibration_date = "2008-02-11" ;
		tsg:intake_depth = "4 ft" ;
		tsg:pipe_length_from_external_water_to_thermosalinograph_meters = "1.1" ;
		tsg:temp_coefficient_G = "4.12651 e -3" ;
		tsg:temp_coefficient_H = "5.84245 e -4" ;
		tsg:temp_coefficient_I = "1.70768 e -6" ;
		tsg:temp_coefficient_J = "-2.49174 e -6" ;
		tsg:temp_coefficient_F0 = "1000.0" ;
		tsg:cond_coefficient_G = "-4.08750" ;
		tsg:cond_coefficient_H = "4.87380 e -1" ;
		tsg:cond_coefficient_I = "1.35767 e -3" ;
		tsg:cond_coefficient_J = "-3.70493 e -5" ;
		tsg:cond_coefficient_CPcor = "-9.5700 e -8" ;
		tsg:cond_coefficient_CTcor = "3.2500 e -6" ;
	byte tmsr(trajectory) ;
		tmsr:long_name = "hull mounted thermistor at thermosalinograph intake" ;
		tmsr:nodc_name = "thermistor" ;
		tmsr:make_model = "n/a" ;
		tmsr:serial_number = "n/a" ;
		tmsr:intake_depth_meters = "n/a" ;
		tmsr:calibration_date = "n/a" ;
		tmsr:temp_coefficient_A0 = "n/a" ;
		tmsr:temp_coefficient_A1 = "n/a" ;
		tmsr:temp_coefficient_A2 = "n/a" ;
		tmsr:temp_coefficient_A3 = "n/a" ;
		tmsr:temp_slope = "n/a" ;
		tmsr:temp_offset = "n/a" ;
	byte sstr(trajectory) ;
		sstr:long_name = "hull mounted thermistor at sea surface" ;
		sstr:nodc_name = "thermistor" ;
		sstr:make_model = "n/a" ;
		sstr:serial_number = "n/a" ;
		sstr:depth_meters = "n/a" ;
		sstr:calibration_date = "n/a" ;
	byte flag_a(trajectory, obs) ;
		flag_a:long_name = "QC flag-platform identification" ;
		flag_a:flag_values = 0b, 1b ;
		flag_a:flag_meanings = "fail pass" ;
		flag_a:comment = "The platform must have a valid call sign" ;
		flag_a:coordinates = "time lat lon" ;
		flag_a:grid_mapping = "crs" ;
	byte flag_b(trajectory, obs) ;
		flag_b:long_name = "QC flag-impossible date" ;
		flag_b:flag_values = 0b, 1b ;
		flag_b:flag_meanings = "fail pass" ;
		flag_b:comment = "The date and time of an observation have to be correct. Valid 4 digit year, month range of 1 to 12, day range for corresponding month, and that the hour-minute-seconds are in the correct ranges" ;
		flag_b:coordinates = "time lat lon" ;
		flag_b:grid_mapping = "crs" ;
	byte flag_c(trajectory, obs) ;
		flag_c:long_name = "QC flag-impossible location" ;
		flag_c:flag_values = 0b, 1b ;
		flag_c:flag_meanings = "fail pass" ;
		flag_c:comment = "This test requires correct latitude and longitude values for the observations. Latitude within the range -90 to 90 and longitude within the range -180 to 180." ;
		flag_c:coordinates = "time lat lon" ;
		flag_c:grid_mapping = "crs" ;
	byte flag_d(trajectory, obs) ;
		flag_d:long_name = "QC flag-position on land step" ;
		flag_d:flag_values = 0b, 1b ;
		flag_d:flag_meanings = "fail pass" ;
		flag_d:comment = "This test requires that the latitude and longitude of the observation is located at sea. The ETOPO2/TerrainBase file is used to see if each data point is located at sea." ;
		flag_d:coordinates = "time lat lon" ;
		flag_d:grid_mapping = "crs" ;
	byte flag_e(trajectory, obs) ;
		flag_e:long_name = "QC flag-impossible speed" ;
		flag_e:flag_values = 0b, 1b ;
		flag_e:flag_meanings = "fail pass" ;
		flag_e:comment = "The speed between 2 observations cannot exceed a maximum value. If the speed is higher than permitted for the platform (usually cargo or research ship), the location, date or identification of the platform may be incorrect. The speed is calculated between an observation and the previous one. If there is no previous observation, the test is correct." ;
		flag_e:coordinates = "time lat lon" ;
		flag_e:grid_mapping = "crs" ;
	byte flag_f(trajectory, obs) ;
		flag_f:long_name = "QC flag-global ranges" ;
		flag_f:flag_values = 0b, 1b ;
		flag_f:flag_meanings = "temp_or_sal_not_within_valid_global_ranges temp_or_sal_within_valid_global_ranges" ;
		flag_f:comment = "This test applies a gross filter on observed values for temperature and salinity. It needs to accommodate all of the expected extremes encountered in the oceans. The temperature within range -2.5 to 45.0 degree Celsius and salinity within range 0.0 to 60 PSU" ;
		flag_f:coordinates = "time lat lon" ;
		flag_f:grid_mapping = "crs" ;
	byte flag_g(trajectory, obs) ;
		flag_g:long_name = "QC flag-regional ranges" ;
		flag_g:flag_values = 0b, 1b ;
		flag_g:flag_meanings = "temp_or_sal_not_within_valid_global_ranges temp_or_sal_within_valid_global_ranges" ;
		flag_g:comment = "The test applies to only certain regions of the workd, where conditions can be further qualified, For example, specific ranges for observations from the Mediterranean and Red Seas further restrict what are considered sensible values.  The Red Sea is defined by the region (10N 40E), (20N 50E), (30N 30E), (10N 40E), and the Mediterranean Sea by the region (30N 6W), (30N 40E), (40N 35E), (42N 20E), (50N 15E), (40N 5E), (30N 6W). For the Red Sea, temperature within range 21.7 to 40.0 degree Celsius and salinity within range 0.0 to 41.0 PSU. For the Mediterranean Sea, temperature within range 10.0 to 40.0 degree Celsius and salinity within range 0.0 to 40.0 PSU" ;
		flag_g:coordinates = "time lat lon" ;
		flag_g:grid_mapping = "crs" ;
	byte flag_h(trajectory, obs) ;
		flag_h:long_name = "QC flag-spike test" ;
		flag_h:flag_values = 0b, 1b ;
		flag_h:flag_meanings = "temp_or_sal_failed_spike_test temp_or_sal_passed_spike_test" ;
		flag_h:comment = "The difference between sequential measurements, where one measurement is quite different than adjacent ones, is a spike in both size and gradient. Test value= |V2-(V3+V1)/2| - |(V3-V1)/2|, where V2 is the measurement being tested as a spike, and V1 and V3 are the previous and next. For temperature, the V2 value is flagged as wrong when the test value exceeds 6.0 degree Celsius. For salinity, the V2 value is flagged as wrong when the test value exceeds 0.9 PSU." ;
		flag_h:coordinates = "time lat lon" ;
		flag_h:grid_mapping = "crs" ;
	byte flag_i(trajectory, obs) ;
		flag_i:long_name = "QC flag-constant value" ;
		flag_i:flag_values = 0b, 1b ;
		flag_i:flag_meanings = "value_constant value_not_constant" ;
		flag_i:comment = "The test is failed when there is no difference in the values of the measured parameters during a six hour period." ;
		flag_i:coordinates = "time lat lon" ;
		flag_i:grid_mapping = "crs" ;
	byte flag_j(trajectory, obs) ;
		flag_j:long_name = "QC flag-gradient test" ;
		flag_j:flag_values = 0b, 1b ;
		flag_j:flag_meanings = "fail pass" ;
		flag_j:comment = "The test is failed when the difference between adjacent measurements is too steep. Test value = |V2-(V3+V1)/2|, where V2 is the measurement being tested as a spike, and V1 and V3 are the previous and next values. For water temperature, the V2 value is flagged as wrong when the test value exceeds 9.0 degree Celsius. For salinity, the V2 value is flagged as wrong when the test value exceeds 1.5." ;
		flag_j:coordinates = "time lat lon" ;
		flag_j:grid_mapping = "crs" ;
	byte flag_k(trajectory, obs) ;
		flag_k:long_name = "QC flag-climatology and NCEP weekly analysis" ;
		flag_k:flag_values = 0b, 1b ;
		flag_k:flag_meanings = "fails_climatology passes_climatology" ;
		flag_k:comment = "Each measurement is compared against a monthly climatology (Levitus 2001, 1 degree by 1 degree, monthly) and against the NCEP weekly analysis fields. The test fails if |V1-V2|>3*Sigma, where V1 is the value to be controlled, V2 is the value of the climatology or NCEP field, and Sigma is the standard deviation of the climatology." ;
		flag_k:coordinates = "time lat lon" ;
		flag_k:grid_mapping = "crs" ;
	byte flag_l(trajectory, obs) ;
		flag_l:long_name = "QC flag-buddy check" ;
		flag_l:flag_values = 0b, 1b ;
		flag_l:flag_meanings = "fails_buddy_check passes_buddy_check" ;
		flag_l:comment = "Each measurement is compared with profiling floats, XBTs, CTDs, thermistor chain, and drifter data (referred here as buddy) within 100 km and plus/minus 5 days of the TSG measurement. Test value = |V1-V2|, where V1 is the value to be controlled and V2 is the value of the buddy. For temperature, the V1 value is flagged when the test value exceeds 0.5 degree Celsius. For salinity, the V1 value is flagged when the test value exceeds 0.2 PSU." ;
		flag_l:coordinates = "time lat lon" ;
		flag_l:grid_mapping = "crs" ;
	byte crs(trajectory) ;
		crs:grid_mapping_name = "latitude_longitude" ;
		crs:epsg_code = "EPSG:4326" ;
		crs:longitude_of_prime_meridian = 0. ;
		crs:semi_major_axis = 6378137. ;
		crs:inverse_flattening = 298.257223563 ;

// global attributes:
		:title = "Underway sea surface temperature and salinity aboard the David Starr Jordan on 20080615." ;
		:summary = "The data being submitted to NODC contain information about temperature and salinity obtained with the use of thermosalinographs (TSG) installed in ships of the NOAA fleet and other cargo and cruise ships. The data is transmitted to AOML/NOAA in real-time and submitted to a quality control procedure developed at AOML based on the Global Ocean Surface Underway Data Pilot Project (GOSUD) real-time control test. Data approved in these tests are submitted to the GTS. The data set submitted to NODC for distribution constitute the complete data set received by AOML with the corresponding flags after the quality control." ;
		:institution = "US DOC; NOAA; Office of Marine and Aviation Operations" ;
		:source = "insitu observation" ;
		:uuid = "73d10173-333b-4525-af74-523c451c56e2\n",
			"" ;
		:id = "AOML-TSG_WTDK_20080615" ;
		:naming_authority = "gov.noaa.aoml.phod" ;
		:references = "http://www.aoml.noaa.gov/phod/tsg/index.php" ;
		:platform = "plt" ;
		:geospatial_lat_min = 33.29583 ;
		:geospatial_lat_max = 34.338 ;
		:geospatial_lon_min = -120.77133 ;
		:geospatial_lon_max = -119.6485 ;
		:geospatial_lat_units = "degrees_north" ;
		:geospatial_lon_units = "degrees_east" ;
		:time_coverage_start = "2008-06-15T00:00:19Z" ;
		:time_coverage_end = "2008-06-15T23:59:49Z" ;
		:date_created = "2011-10-25T22:24:14Z" ;
		:creator_name = "US DOC; NOAA; NESDIS; National Oceanographic Data Center" ;
		:creator_url = "http://www.nodc.noaa.gov" ;
		:creator_email = "NODC.Services@noaa.gov" ;
		:project = "AOML-TSG" ;
		:processing_level = "Synthesized Products" ;
		:featureType = "trajectory" ;
		:cdm_data_type = "Trajectory" ;
		:Conventions = "CF-1.6" ;
		:Metadata_Conventions = "Unidata Dataset Discovery v1.0" ;
		:standard_name_vocabulary = "NetCDF Climate and Forecast (CF) Metadata Convention Standard Name Table v23" ;
		:keywords_vocabulary = "GCMD Science Keywords" ;
		:keywords = "Oceans > Ocean Temperature > Water Temperature, Oceans > Salinity/Density > Conductivity, Oceans > Salinity/Density > Salinity" ;
		:comment = "NOAA/AOML/PhOD assessed the quality of the data using an automated quality control flagging procedure." ;
		:history = "This netCDF file was created by the National Oceanographic Data Center using the original file from the ship and the corresponding quality controlled file created by AOML." ;
		:nodc_template_version = "NODC_Trajectory_Template_v1.1" ;
}

netcdf \00000110200000-NODC-L4_GHRSST-SSTskin-AVHRR_Pathfinder-PFV5.0_Daily_Climatology_1982_2008_DayNightCombined-v02.0-fv01.0 {
dimensions:
	lat = 4096 ;
	lon = 8192 ;
	nv = 2 ;
	time = 1 ;
variables:
	int time(time) ;
		time:standard_name = "time" ;
		time:long_name = "reference time of climatological sst field" ;
		time:climatology = "climatology_bounds" ;
		time:units = "seconds since 1981-01-01 00:00:00" ;
		time:axis = "T" ;
		time:calendar = "Gregorian" ;
	int climatology_bounds(time, nv) ;
		climatology_bounds:units = "seconds since 1981-01-01 00:00:00" ;
		climatology_bounds:comment = "This variable defines the bounds of the climatological time period in this file. It contains two time elements: the first specifies the beginning of the first subinterval (in this case, one day); the second specifies the end of the last subinterval used to evaluate the daily climatological SST for this file." ;
	float lat(lat) ;
		lat:standard_name = "latitude" ;
		lat:units = "degrees_north" ;
		lat:valid_min = -90.f ;
		lat:valid_max = 90.f ;
		lat:axis = "Y" ;
		lat:bounds = "lat_bounds" ;
	float lat_bounds(lat, nv) ;
		lat_bounds:units = "degrees_north" ;
		lat_bounds:comment = "This variable defines the latitude values at the north and south bounds of every 4km pixel." ;
	float lon(lon) ;
		lon:standard_name = "longitude" ;
		lon:units = "degrees_east" ;
		lon:valid_min = -180.f ;
		lon:valid_max = 180.f ;
		lon:axis = "X" ;
		lon:bounds = "lon_bounds" ;
	float lon_bounds(lon, nv) ;
		lon_bounds:units = "degrees_east" ;
		lon_bounds:comment = "This variable defines the longitude values at the west and east bounds of every 4km pixel." ;
	byte crs(time) ;
		crs:_Unsigned = "true" ;
		crs:grid_mapping_name = "latitude_longitude" ;
		crs:longitude_of_prime_meridian = 0. ;
		crs:semi_major_axis = 6378137. ;
		crs:inverse_flattening = 298.257223563 ;
		crs:comment = "This is a container variable that describes the grid_mapping used by the data in this file. This variable does not contain any data; only information about the geographic coordinate system." ;
	short analysed_sst(time, lat, lon) ;
		analysed_sst:_CoordinateAxes = "time lat lon " ;
		analysed_sst:standard_name = "sea_surface_skin_temperature" ;
		analysed_sst:long_name = "analysed climatological sea surface temperature" ;
		analysed_sst:cell_methods = "time: mean within years time: mean over years" ;
		analysed_sst:units = "kelvin" ;
		analysed_sst:add_offset = 273.15 ;
		analysed_sst:scale_factor = 0.01 ;
		analysed_sst:valid_min = -180s ;
		analysed_sst:valid_max = 4500s ;
		analysed_sst:_FillValue = -32768s ;
		analysed_sst:grid_mapping = "crs" ;
		analysed_sst:ancillary_variables = "analysis_error sea_ice_fraction mask" ;
		analysed_sst:comment = "Daily climatological skin temperature of the ocean, derived from harmonic analysis of the AVHRR Pathfinder Version 5.0 sea surface temperature time series from 1982-2008." ;
	short analysis_error(time, lat, lon) ;
		analysis_error:_CoordinateAxes = "time lat lon " ;
		analysis_error:standard_name = "sea_surface_temperature_error" ;
		analysis_error:long_name = "estimated error standard deviation of climatological SST" ;
		analysis_error:cell_methods = "time: mean within years time: mean over years" ;
		analysis_error:units = "kelvin" ;
		analysis_error:add_offset = 0. ;
		analysis_error:scale_factor = 0.01 ;
		analysis_error:valid_min = 0s ;
		analysis_error:valid_max = 32767s ;
		analysis_error:_FillValue = -32768s ;
		analysis_error:grid_mapping = "crs" ;
		analysis_error:comment = "This field is taken from the standard deviation maps generated during calculation of the \"classic,\" or mean, daily climatology for Pathfinder Version 5.0. The original layers can be found at http://data.nodc.noaa.gov/opendap/pathfinder/Version5.0_CloudScreened/Daily/FullRes/climatology/contents.html in the ClimSTDV7_daynitavg layer." ;
	byte sea_ice_fraction(time, lat, lon) ;
		sea_ice_fraction:_Unsigned = "true" ;
		sea_ice_fraction:_CoordinateAxes = "time lat lon " ;
		sea_ice_fraction:standard_name = "sea_ice_area_fraction" ;
		sea_ice_fraction:long_name = "climatological sea ice area fraction" ;
		sea_ice_fraction:cell_methods = "time: mean over years" ;
		sea_ice_fraction:units = "1" ;
		sea_ice_fraction:add_offset = 0. ;
		sea_ice_fraction:scale_factor = 0.01 ;
		sea_ice_fraction:valid_min = 0b ;
		sea_ice_fraction:valid_max = 100b ;
		sea_ice_fraction:_FillValue = -128b ;
		sea_ice_fraction:grid_mapping = "crs" ;
		sea_ice_fraction:ancillary_variables = "sea_ice_fraction_error" ;
		sea_ice_fraction:source = "EUMETSAT OSISAF Global Daily Sea Ice Concentration Reprocessing Data Set" ;
		sea_ice_fraction:comment = "Sea ice concentration data were taken from the EUMETSAT Ocean and Sea Ice Satellite Application Facility (OSISAF) Global Daily Sea Ice Concentration Reprocessing Data Set (http://accession.nodc.noaa.gov/0068294). The data were reprojected and interpolated from their original polar stereographic projection at 10km spatial resolution to the 4km Pathfinder Version 5.0 grid. A classic daily mean climatology was then calculated." ;
	byte sea_ice_fraction_error(time, lat, lon) ;
		sea_ice_fraction_error:_Unsigned = "true" ;
		sea_ice_fraction_error:_CoordinateAxes = "time lat lon " ;
		sea_ice_fraction_error:long_name = "standard deviation of climatological sea ice area fraction" ;
		sea_ice_fraction_error:cell_methods = "time: mean over years" ;
		sea_ice_fraction_error:units = "1" ;
		sea_ice_fraction_error:add_offset = 0. ;
		sea_ice_fraction_error:scale_factor = 0.01 ;
		sea_ice_fraction_error:valid_min = 0b ;
		sea_ice_fraction_error:valid_max = 100b ;
		sea_ice_fraction_error:_FillValue = -128b ;
		sea_ice_fraction_error:source = "EUMETSAT OSISAF Global Daily Sea Ice Concentration Reprocessing Data Set" ;
	byte mask(time, lat, lon) ;
		mask:_Unsigned = "true" ;
		mask:_CoordinateAxes = "time lat lon " ;
		mask:long_name = "land sea ice lake bit mask" ;
		mask:valid_min = 0b ;
		mask:valid_max = 8b ;
		mask:flag_meanings = "ocean land lake_surface sea_ice river_surface" ;
		mask:flag_values = 0b, 1b, 2b, 4b, 8b ;
		mask:grid_mapping = "crs" ;
		mask:source = "Land pixels were determined by rasterizing to 4km the Global Self-consistent Hierarchical High-resolution Shoreline (GSHHS) Database from the NOAA National Geophysical Data Center using a 50 percent area threshold. Inland water bodies (rivers and lakes) were determined by rasterizing to 4km the US World Wildlife Fund Global Lakes and Wetlands Database using a 50 percent area threshold." ;

// global attributes:
		:Conventions = "CF-1.6" ;
		:title = "AVHRR Pathfinder Version 5.0 and 5.1 Harmonic Climatology for Daily Day/Night Combined Sea Surface Temperature, 1982-2008" ;
		:summary = "This netCDF-4 file contains global 4km daily day/night combined sea surface temperature climatology values for yearday 010 (Jan 10) derived from harmonic fit analysis of 5-day averaged AVHRR Pathfinder Version 5.0/5.1 sea surface temperature data for 1982-2008." ;
		:references = "http://pathfinder.nodc.noaa.gov and Casey, K.S., T.B. Brandon, P. Cornillon, and R. Evans: The Past, Present and Future of the AVHRR Pathfinder SST Program, in Oceanography from Space: Revisited, eds. V. Barale, J.F.R. Gower, and L. Alberotanza, Springer, 2010. DOI: 10.1007/978-90-481-8681-5_16." ;
                :featureType = "grid" ;
                :cdm_data_type = "Grid" ;
		:institution = "NODC" ;
		:history = "compute_harmonic_clim_col.m, compute_climatology.m" ;
		:comment = "AVHRR Pathfinder data of quality flag 7 only" ;
		:license = "These data are available for use without restriction." ;
		:id = "AVHRR_Pathfinder-NODC-L4-DailyClimatology-v5.0" ;
		:naming_authority = "org.ghrsst" ;
		:product_version = "PFV5.0 and PFV5.1" ;
		:netcdf_version_id = "4.1.2" ;
		:gds_version_id = "2.0" ;
		:file_quality_level = 3. ;
		:source = "AVHRR Pathfinder Version 5.0 and 5.1 5-day day/night combined SST, Quality flag 7 only" ;
		:platform = "NOAA-07, NOAA-09, NOAA-11, NOAA-14, NOAA-16, NOAA-17, NOAA-18" ;
		:sensor = "AVHRR_GAC" ;
		:Metadata_Conventions = "Unidata Dataset Discovery v1.0" ;
                :nodc_template_version = "NODC_NetCDF_Grid_Template_v1.1" ;
		:metadata_link = "http://accession.nodc.noaa.gov/0071181" ;
		:standard_name_vocabulary = "NetCDF Climate and Forecast (CF) Metadata Convention Standard Name Table v23" ;
		:westernmost_longitude = -180.f ;
		:easternmost_longitude = 180.f ;
		:southernmost_latitude = -90.f ;
		:northernmost_latitude = 90.f ;
		:spatial_resolution = 0.0439 ;
		:geospatial_lat_units = "degrees_north" ;
		:geospatial_lat_resolution = 0.0439 ;
		:geospatial_lon_units = "degrees_east" ;
		:geospatial_lon_resolution = 0.0439 ;
		:geospatial_lon_min = -180.f ;
		:geospatial_lon_max = 180.f ;
		:geospatial_lat_min = -90.f ;
		:geospatial_lat_max = 90.f ;
		:geospatial_vertical_min = 0.f ;
		:geospatial_vertical_max = 0.f ;
		:geospatial_vertical_units = "m" ;
		:geospatial_vertical_resolution = "point" ;
		:geospatial_vertical_positive = "down" ;
		:acknowledgment = "Please acknowledge the use of these data with the following statement: These data were provided by GHRSST and the US National Oceanographic Data Center." ;
		:creator_name = "Kenneth S. Casey" ;
		:creator_email = "Kenneth.Casey@noaa.gov" ;
		:creator_url = "http://pathfinder.nodc.noaa.gov" ;
		:project = "Group for High Resolution Sea Surface Temperature, Pathfinder" ;
		:publisher_name = "GHRSST Project Office" ;
		:publisher_email = "ghrsst-po@nceo.ac.uk" ;
		:publisher_url = "http://www.ghrsst.org" ;
		:contributor_name = "Robert Evans" ;
		:contributor_role = "scienceParty" ;
		:processing_level = "L4" ;
		:cdm_data_type = "Grid" ;
		:keywords = "Oceans > Ocean Temperature > Sea Surface Temperature" ;
		:keywords_vocabulary = "NASA Global Change Master Directory (GCMD) Science Keywords" ;
		:date_created = "20110811T194351Z" ;
		:date_modified = "20110811T194351Z" ;
		:date_issued = "20110822T090000Z" ;
		:start_time = "00000110T080000Z" ;
		:time_coverage_start = "00000110T080000Z" ;
		:stop_time = "00000111T075959Z" ;
		:time_coverage_end = "00000111T075959Z" ;
		:time_coverage_resolution = "P1D" ;
		:time_coverage_duration = "P1D" ;
		:uuid = "4b066e2a-b791-42ea-94b6-828c1b2b24fe" ;
}

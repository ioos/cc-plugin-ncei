netcdf NCEI_TimeSeries_Orthogonal {
dimensions:
       time = 1;
variables:
        double time(time) ;
                time:long_name = "Time" ; 
                time:standard_name = "time" ; 
                time:units = "seconds since 1970-01-01 00:00:00 0:00" ; 
                time:calendar = "gregorian" ; 
                time:axis = "T" ; 
                time:ancillary_variables = "" ; 
                time:comment = "Time" ; 
        float lat ;
                lat:long_name = "Latitude" ; 
                lat:standard_name = "latitude" ; 
                lat:units = "degrees_north" ; 
                lat:axis = "Y" ; 
                lat:valid_min = -90.0f ; 
                lat:valid_max = 90.0f ; 
                lat:_FillValue = -9999.0f;
                lat:ancillary_variables = "" ; 
                lat:comment = "" ; 
       float lon ; 
                lon:long_name = "Longitude" ; 
                lon:standard_name = "longitude" ; 
                lon:units = "degrees_east" ; 
                lon:axis = "X" ; 
                lon:valid_min = -180.0f ; 
                lon:valid_max = 180.0f ; 
                lon:_FillValue = -9999.0f;
                lon:ancillary_variables = "" ; 
                lon:comment = "" ; 
        float z ;
                z:long_name = "Depth Below Sea Surface" ; 
                z:standard_name = "depth" ; 
                z:units = "m" ; 
                z:axis = "Z" ; 
                z:positive = "down" ; 
                z:valid_min = 0.0f ; 
                z:valid_max = 1000.0f ; 
                z:_FillValue = -9999.0f;
                z:ancillary_variables = "" ; 
                z:comment = "" ; 

        float temperature(time) ;
                temperature:long_name = "Sea Water Temperature" ; 
                temperature:standard_name = "sea_water_temperature" ; 
                temperature:ncei_name = "" ; 
                temperature:units = "" ; 
                temperature:scale_factor = 0.0f ; 
                temperature:add_offset = 0.0f ; 
                temperature:_FillValue = 0.0f ; 
                temperature:missing_value = 0.0f ; 
                temperature:valid_min = 0.0f ; 
                temperature:valid_max = 0.0f ; 
                temperature:coordinates = "time lat lon z" ; 
                temperature:coverage_content_type = "" ; 
                temperature:grid_mapping = "crs" ; 
                temperature:source = "" ; 
                temperature:references = "" ; 
                temperature: cell_methods = "" ; 
                temperature:ancillary_variables = "temperature_qc" ; 
                temperature:platform = "platform_id" ; 
                temperature:instrument = "instrument_id";
                temperature:comment = "" ; 

        int temperature_qc(time);  
                temperature_qc:standard_name= "" ; 
                temperature_qc:long_name = "" ; 
                temperature_qc:flag_values = ""; 
                temperature_qc:flag_meanings = "" ; 
                temperature_qc:references = "" ; 
                temperature_qc:comment = "" ; 

        int platform_id; 
                platform_id:long_name = "" ; 
                platform_id:comment = "" ; 
                platform_id:call_sign = "" ; 
                platform_id:ncei_code = ""; 
                platform_id:wmo_code = "";
                platform_id:imo_code  = "";

        int instrument_id; 
                instrument_id:long_name = "" ; 
                instrument_id:comment = "" ; 
        double crs; 
                crs:grid_mapping_name = "latitude_longitude"; 
                crs:epsg_code = "EPSG:4326" ; 
                crs:semi_major_axis = 6378137.0d ; 
                crs:inverse_flattening = 298.257223563d ; 



       :ncei_template_version = "NCEI_NetCDF_TimeSeries_Orthogonal_Template_v2.0" ; 
       :featureType = "timeSeries" ; 
       :title = "Example Time Series Dataset" ; 
       :summary = "This dataset is just for demonstration and testing purposes" ; 
       :keywords = "examples" ; 
       :Conventions = "CF-1.6" ; 
       :id = "some-uuid" ; 
       :naming_authority = "com.asascience" ; 
       :history = "Generated for testing purposes" ; 
       :source = "Luke's brain" ; 
       :processing_level = "raw" ; 
       :comment = "Just for testing purposes" ; 
       :acknowledgment = "I'd like to thank the academy" ; 
       :license = "freely distributable but for testing only" ; 
       :standard_name_vocabulary = "NetCDF Climate and Forecast (CF) Metadata Convention Standard Name Table \"29\"" ; 
       :Metadata_Conventions = "Unidata Dataset Discovery v1.0"
       :date_created = "2016-05-20" ; 
       :creator_name = "Luke Campbell" ; 
       :creator_email = "omitted" ; 
       :creator_url = "https://github.com/ioos/compliance-checker/" ; 
       :institution = "RPS ASA" ; 
       :project = "IOOS Compliance Checker" ; 
       :publisher_name = "Luke Campbell" ; 
       :publisher_email = "omitted" ; 
       :publisher_url = "https://github.com/ioos/compliance-checker/" ; 
       :geospatial_lat_min = 0.0f ; 
       :geospatial_lat_max = 0.0f ; 
       :geospatial_lon_min = 0.0f ; 
       :geospatial_lon_max = 0.0f ; 
       :geospatial_vertical_min = 0.0f ; 
       :geospatial_vertical_max = 0.0f ; 
       :geospatial_vertical_positive = "down" ; 
       :time_coverage_start = "2016-05-17T00:00:00Z" ; 
       :time_coverage_end = "2016-05-18T00:00:00Z" ; 
       :time_coverage_duration = "P1D" ; 
       :time_coverage_resolution = "point" ; 
       :uuid = "another-uuid" ; 
       :sea_name = "Mid-Atlantic Bight" ; 
       :contributor_name = "Luke Campbell" ; 
       :contributor_role = "Owner" ; 
       :geospatial_lat_units = "degrees_north" ; 
       :geospatial_lon_units = "degrees_east"; 
       :geospatial_vertical_units = "m" ; 
       :date_modified = "2016-05-20" ; 
       :keywords_vocabulary = "" ; 
       :platform = "" ; 
       :instrument = "instrument_id" ; 
       :cdm_data_type = "Station" ; 
       :metadata_link = "http://google.com/" ; 
       :references = "http://google.com/" ; 
       
      
}
